`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WXMgGoH0V1HcubY4hXKMghp9Z8XrMh09TFuiMytgMPlB3bDvsBffXlJu0elhS5XNp2rkE45zzIER
kLqAza7KTA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Zir/Ug+A/WnX12oS0+9Inww916NGKNU9LAmTuV0QareNJzykYy0GM/uDdWuRnBSkkPRUv8muQwqu
uryEkLvLO3o9QfjC9jrEWz2Ep83oQaPOVySRRsFplMq2seM9gnQNpKyBYWRLmi1y3LiVJCyudlij
FbYZiN832GgcveDITos=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qSmSI2AzVfH0PCcOA7lDlP82yNQSNwIcoYI4D1QLyxCjx3qLvbI6tlO9AoVNQ5nhlnG558/dyvvE
AcqaZEIoDtjt6JbNzI4utc8xEB+6NKsHbmQn5uJg02u8qyKXrid7zvYuSb/rEM+aRkE5HeTqQm5E
dIkRAmYuACagsEHug38qprbo50TCN+ilsyNr3964QZEkSTGtCVqKa1f66jrBWj/n7nliqe2Lpinl
+u0Z1UPYB0HAzDYF15gB3ZsIFcsm4xyaBbzLoDDFCQXF/Oi2IXrUn3QeOUr6EVpbInAjDY3eKKTc
/jmi9bf3rflmaMO+hJ6WY37q4mVK6Ik9FACTvA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Hu1g7ldnrGKXqJ3jd2VNpp7RS6+QnqBCUvcj788HuY/zbGCh2psBSwEYarHM4SRGyPIxKuyNNNSU
v8lKHJH/cI+eYKV68+L+9ie7CwQ/uz1JrD1Ow57FuJM4WTqnaoBUw8ljgXmb43UZiRtDrhxeiNGw
aVK81eyeRLEIiNG/9Qo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fz0NxXH4fercPobk/9V/c3BsrWVixhUxSd80FE8LZJd6zUx5YzGyQnwQB6BtvzKWMfsORfdRfaSg
Xmw4YxiV7AyKpKQtW5lT/Vmac9k9RVwGkmcLkxC1bhcj4DbZ7HUfEgnglSPPmktjDBjqHAgBZQXW
qxjMkZsM3zgZJ6zpI7N4zo+4bzhoz4xQZjKP+2XUA+epHj+SD/4HrTkLRyd6Ahk2IqQW9N2IEynP
MPKGsRv6O+AwL+Lqgknd/v/hTY3ZE5YffjWHfepoqVVxBbY9ulUmnAmtMNQye7i80ZfAPs/18xUY
MDx8O6LSRKMO4s5U63EfUyEsO2u1KMudT83uVw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10432)
`protect data_block
wW8P7V+nTkMAaoGxyhyUNIi6DaKGpq2ZoJ4jNSZG+s8ISWYTSSp7B5wQd2zGZhrg/LZnN/s2ohoa
KJfxk3w2oAO7FNDzZnuVZPuq9B3vQWc8fORAH7s9zMJaYjh6Jvxu7RfxY3y2jARGJ2L56iVZhABG
3cHygOrsbE8expIrIhIYYzvqPBgW18ytD0g3+vphu1Tu07iYQ92X9ewJeEhB7PqU3UttMbCLnvUr
kNMv52qYT+W4Qvic8gog5UaQ6ZxxHQFJnGAI+6St0Crxpb9wIcoXK8YOBDGrjrLh2DtIpK+rPrJw
mpmN7+frHUr5skOU95zcOlxGb2YfZ6ZR7z8J4SN8FIoWns4f3WSWHJllB5FHyaZz5dR3RGaysbGX
7NMgQe8vNOBcnBu5iD/XTs8nHgoNgkhkgs6ynkUc3u2ZfG07t7bCEIRgiLwmSv3xiD2FKxL9BGjG
CYr2EYmcP6zGOUWrnuH/DLIINXTm8w99Jl5ULENR63KGQQAbfNT3zX/BW34tWrgxRRUJn2jmattw
fo97ezft/iktVw8jwEX8gpSB64BLkXQyM6aVCBKm4OgrGm3iV08vKF9j1QImLWcB0pfJ5W4ea3m3
SGLhmCI5cnrV/fUUi1GCGGGi++e88GBLEbD+VTUSNftx9LH6YQoL9A9UDMOIkX484mqQ6F2bux7W
JeImvovwUs3Z+UHzn9ZP+KmV1PVQbC41ET+sjB2Snll/uk0JhN3CQ0z5Ih1IsBrDRzUVPi2PlXjj
+5vwuIzYopnAh0CGLFYZsz9OjuFnGWVh6VnotdAx98hpHVf1hQqZrJYQRQ6miI9Et1+VRMd5pxg8
BFj/cnOdkSYVz4zKjQdB55UaYVzBAUdibWVJFWQd36ANzV+SV7zbX2AJP86ESWbvD6eCqJ12ZciJ
N1/ZcB7dSgnNjcXIm0gRK1VtHIjBejE/GLnxIE0jgcG1cKUVCOuuaEZsczf8mYNDIOQkXoNbkfZT
GLxI2nuVUST87+3AyB578FTA/WcHEn36+Q8g+IJvzEc/AtI/0xRDYn5pHVqTDUT99logVOacW/sN
O8CYp2CD2fh2+GtavTFWYlefWNGQ5WhaiVYlzZjzJVUa0FDAfwjNfsZIJGDueOcDGSeqY6VJDHtJ
94+m9jB3Ikgo5mopiCgJKt5Hpl3FIiFgbu5yXEr282QGbCrKqiSAahXyCdJNc0deZaih6hQE7Hpi
9ICriabFPGbuU3AWioPGNzNdKtELlkW4CPvVAbIe24RtN8uPyGdUVfhnknVCMPWSDII5LakyffNi
zVUCtFCfo1bLVoFdJSADHUq/sQ83nlBWP+fTeE7UtrVM4REJLSKBs/wtU0XaSxWkXUzppFb+dNv3
FOmSppWqyMkbE36lRbT4062DSVMemFphTve7sOi56jehOpbudi3XUfEJWWPAuZnJTNAY7ilfQbqY
IDnAb2yiZqGpsA3mh2OOLj8GgzAWNyVJ1nRtnN87vWlNk3P8osZlUhKvCziVdmXtXJ3G5L33djp0
XImzO3/BIegsLKVvKxkYteFeruZm5P+Hb1IV4gnTR7Q/KrOcNyn8tDsBgDQAUWVThdGx50bWomV7
hqLcpinqR21DpUmPsW3WZe/Fn27CI7JtJdp1AQOS+9c28TukNeuCtVKoplgW+MGUIAq1AwZfDclo
fJ3whfiy7/hu1xsu+eHBt2XD26v84g9OpY0Rm0jlWM9EinjJ+PugaqSl93G/VhKISIJ8xGsNLPYn
GqD8UfYRcMrt8315kRVNR0AqGhZ8h3GqYNCsEqUAlZkF9esDO9XQVALmI5Nemrpw0n9oHHze/6lO
tAkVzGvHSyG37cSkveyz233N60mWEAZHW59zYUM8o94p422yZdSgHwjbZ3aDnEktWCUUXpfF+yKR
dhaVbUc2QmjusBHojoBOFT4deNr9YVplOrs367pEYctHBEPpWbmg1xXNTNUtbDMZKCfeoAMuYvPh
cMQ1MYGrHppZ5sOdCORDkhuGKQOKY1dOYf0wWHCr39qR8SgJxhm2RJRJqz7uWZrSN5Se7pxLkH6n
84lPuXPpQjCt8KCKUT2GrQwI4wsI5+8IMbzhRQWsLO6kuqxQLJ6F5zgBVDZKhHS+uwQtZi1HojHU
9teQ2hJe+KakbmhdpzN2HWYQjPASrC5+lLkxUJsvl4M1vYLsVAsxOtYXkCLSRVwnjdcEJxbSoxE2
1DXTLGb+T9Tuj/9gsepi8fKD7cKUYM7GrZcdrV1UNM60J3WPuWvlDAMRPhP+pRGdpZ9ZrS7yjQaw
IdgMdxN96vipF5boZ+x1TRzgIQNxjPA/k5C3oHoRSXYvXoUCmKhUFnbNJDWT1LqaBQjQ5Q5v3ext
puOFR33Hm4Yc7PfbayP7mte1I+tgvtO79rpAo+bXHa8gmS2K+Upf5DQqqI7pqZfvV9SSJAhf3aB/
EiFQIvOJslsmbz/OoYbHhM1pIn7lKS0Acb2cy0oxkot/ashFaN515E/atEsromAqB6kaBk+bA7/G
zCKU7v1NBHZPpzdwNhVu74meJ0+OaEjisPOwFXRVSRTJZ18d0CoeCO5eL20C/UJDxm06InoFKjor
pBs5shc88PFRW9V+XJSM+nldKqwzcl+aavgmxPEQgp6VxoDmuutMvHznKp1pGJLw+W4m3SVX9unP
VpIDJHn6rPEg+QP0443/g+T6oUfouDFbiB+2eDWFyXAGmPAl1xGm0Cvl214f6yRySeLJpJozfYZa
UABsnwUWYfnUuhnlmlcLEKm71VCASzumec+l77/c70exJsb9CT93Dr7G4o7R7i4BBC6BsXGF4QLn
H6yEQCmyxKTS9eUytytK4GaBePv8aWzTi0jA+ZLCBHKtpwnKjXi7hL3ct3cGwJIbHH2AlaUYZya+
G7uT9hIY5gh/WIYM9A4VaTP3GLPYQ0Ldxv82SQAsXiCatLW1+uyjvIghh6XMk6GtknCB0/MTJCBV
GmzGB/344bLdz9qUxC9D7z49Ct6yYxyd97pbknB3st0ddtKtY/QEGvJ7y3Iw7g/MUkc2j9Gx8SSc
mPWJfyHEvgeX7dKOgKpcaIu9e/VDJWiSZ5IzXaDSpD0Of26eCGx5tkIG4L9R+5E/AHg3TEtnOdRO
J5xy1L7OrSpaFbC4IUjVVZNTOIancQ3Lwf/qiJ486IMPIGknFXhpHBdFVkHzB7ZD7nuNA1GRQmg+
XcjEoaKEZNNuIOJpJ9HGdRTztK3G14JR5I5p7xw3kxSCpGrva5KCt4rOlyJksOJ3VUpVY3R/a9qj
DHM1z6DMtdCqez9ZhVzYhOYAfNdngIFE0Me+TEi8q06348cyS/CdQufs17xeyolQqhlqE4gpowCu
FJQT8vhM6NLTFSLKYwPS6xR0xwlyiiK7hgT6Axk0rJ2AAeMQVD5MEsJO15kF9U5BGsYGrZz5On6r
C1oVrj5uNQfCYsvEYW1N6BtDxM3ShLNbR5LEgefSqTvIj91bxc8V52YdaY4woWTqx/y6NakRQM1f
keoSTC00mfpurY9YN6Qx7din4G3Uw2aVHV4Wh8IvWF+kUZ+Pie3+fMdnJs/WOvSV2eDJjf5deTab
0C5Dq0BAUqy+i+6cOeaDBuY6rFPDOwDpctAGQuEPofZ8eZR9F2V6Lp6fRGgFmE21pSattpLRs1+m
ySlYOMT2ZAxLi6scdSrylzKg+89CXcV+oxzhL3BgofQOWllNnuPDW40XebGzONlOZwtmcv2NuL0D
K74WB9OoVHFrWmaE3EPZGAwjsurIycAKsNz7K8x4YZRzBPExRUhDw9FF30e2Eo6cMoF5gRP7B+0F
zG+uDU8/gEfgdpd5DnykL0o5QeIdN0TidZOL6CjJmZ5CqXq0nQThuLvC7IQ/8XMApFpdh14PlEBI
3amGDLoT/dpQHFiXLkkjbQirE2PwvTS0JEOIONq4TIk2/ZkJMXfiBUGcyZ9j3gY+1PHO5yjBzql9
rWLx3RuPlWpUnOOPtzzcd2sptpK24DjLuKguZGDH6Zn4fewOSY6yI82fCX553r6whj3OgvI8dkVO
FcGDUnXcVwyIm4uV1Mt62MdJ5lNe+0uK5y23VlRuwggdku/w+EYBYTSj9hgRiCTgVZU7Q5SXnWee
R9Zl7nKlqRTxj8zojvHeHVzwO5Qe/INX2pX9eaUTe0FbwtvskGqUpo5ff3HXN5DFyN2GdKRrQf/c
AQgxS9mSgN8dRQO2Zl6UT9tgAFRe1UTXOmSK2DmOPWjmIirb8cNXzGJHNFNGJ2g4pqqysj9lqy1q
ZTTy0qCaQnhRQhXf+oaXs31kMVrzc9pG5pwCant4rv24yYlmMBoYsn31XsL7LjzwhEjzKiqtL0fg
i76XNFIPg9HJLzKIMdpc6pBcgrILEf01CTGu/pky9EC3Om6MSxx6NWXrFSOVNTsKbvh0WuNUJ4PC
yp9GWxkCdDwayJBV1Txrs+r2MK3h7dTTje2J8qXHq+nm4MV/EpK0i3JwxJzZzBWcyCKHcnNk7ZKF
mNoV0BDJGS8M+kL6nnESaTU56W7OzAjl2lIebY48rRfJ+pHR9B5l9StiAFjCKBf377FSIW0pEIPL
6vwSVYTWla5iyVoqLg3SpB/Qyh30cwNgy5G6kCqvP2sByzEzzzfUIHGGSR6BaqzKUrceKFb2nzEp
+DuKFl7dGM8APiugEmPSXeWFuTAK8OW+62gFprFxxEGcg+1nXnZqPdtrqe+aJsc0Z41mSH9VADMh
kLrkf5MQtYbdgOz5Pt/xhYr5hhZYzaeiltOap3Fezhw++HcdSoQbg4vnWCiE/SouiAl2WSDktzIE
YPmXHXlbwLIITmqRc4/Tj8VjNyIk2GnISxeqAucVvmd9u5rjFpjTS04Z5cDoqzDiQNPKWWdxBprl
h7QZinBc0tsydTOKFU7IcCVYueRcGKAePsp97UyH6/Wx44P4+CIsL7Nozhn8IHk1lwekuTs1w1dU
lEakCSoY42iJfROED871gGDKmJcNjyOV30Fmcy0LQ4+Im8h/SpiZPKPaCzTbIi7aAlqx+OAyluEw
rCn0ouQo4H1sPkgraHvlCrez4THmB16RhdjJpBk3NVeejTkDa4uAoAdCM3nJenHXWhVLGzNK0zOB
bZA6K6yIDb+g+s1p/TxY0h6LwckWOpcfu0buIyFcSwIrJh7vGqsFog0Ybh7i4f6XJoqwEIXwgs4g
pBrXOgcFkI8OIum5giyR8/6LFyhtpoSVV/k2cGniQ5f9vWwD0wDJr9JqmwquKHAeMfqdlUt9sEni
qmmTzk1RAlPw9S1yC6Loink3vCpss26c60635Lwbq6qxAQRJRkwJgRcVKPhlM4FvGmJqQfKzHzOc
7hsG6P//Of7GAcyjI+8YTsJIheVsa7336b5u60n3nHTNTJLuC2ChWUPg1wf6yEfOOH8/OF9UoiHG
3ETavgoxXPdAX7cAA8qPPtCGC7eo0UmUkhKeGxD817ZHo9RgNCYb8lUpNPr3kfJu62lHcJlFDX8x
paEENel58r7SnV+yJxVZTRJ3wPAiMcyRTma1HLSKA2TuRUXmQ9nTYCenCFECHXz4apRbA+crrZsL
swoYY5bivc9FygKZa6x6s5OG4q+x1rciiSuuAOzGukLKjCiyfLlWnCVZqVrLfGmJuoNYXsxRmxBE
86fGPwpFezh6uiEIGd9Dzx6Il7dSr36mrNGZ3dPX0kH82sKHOPa52uGCQp3RsvdPzXJwOGVdLWw5
d3NmHPbayMLnV+uuOI7MXnIlKUL2Re7H5BOkXh9gotuh4dWfn+SyceILWULWie8NHOlP+z6pIfKW
ZMTjoKxYpVZ+vY9w+lzQGXuNBTJqVnr3YL1UaPTgb6uFyAdNTP/h+P6W82VE+/su8Yktw20ydB/G
tvLoqd8ujqcAMhufj+sdLYz4zCl5cntEIKaUK8jzUz2/76mRNkqA8S+88ROXgqZlMobdRbueE9Ly
fwT6T0xnjPIXyZsCsRdVebNrQQWsopYei3KyfElXAgWVCqczP1zfRQpUB3r39rLrRsItQZL77uxt
520ofHACTF/VFnecD1pwYuW9DDdGED79zsvl/1Piwgzh1pU9W9THGYhkBjti/yBeYOcBMrxYvz8D
RegSBjPIQ/U3+5D2HXh486R5zldPxBW0yyQs9FjNYcMKLL70ndruDy6D4rrq1QBgRePOnXgs4H1C
SdPNfNVAFeQf60bQvGKskC1aB6p6c6Q6+ET6s/2Q65vMTowmk4kyigKQOPQbPBh+KRRBI9uXcqTw
A62B/M5nz+8m2gDO5eFPqsOl/YHKnOHBJl+G9lURIbgdUQ6JIgvnDIuATJI1QbpyNUyYIrRVMZxV
ZuyxcDzk3cFU9CPxlmD9n5awPCGc9QrumzXAQ9wwt5vOPESYAJgoc+x78DxDQp2y8wpYyEFJQbWk
EzFTHU6VCfUQweEdWVgmkmn9LY0oV/pa4+S3mnoOnTmyngY9yrqw9OSoKNLFQL33x7D77x3cIYWu
EgjCruCC7Ei1LUpzFrDjkdN6WcDNljUMpFX7nEu5S2HewnjrnhF562j0pubnFbYQU+rBBgdfLDwx
LuPEnfZLB/rGFb6Q67nZMMhJTZsr2NhC80bIHpDZygEXtcE1sbA/IlPpsc/5LT0FXNUMloztYyc9
KFybKbjDDvE4tvU8hCmautIPt2fJOeyvhKY76qP9s/rWOWdZjrG27xNyQPDqYmPZyb7o9fJv1laK
K3ZHhvWnfLaIZxEXZndSYODtNWJ++UTnc/inD4Qf74pXoG3CJPaWXV4X+Y49aVjZuRi399gkqby/
irxQAatploKVdDxR+5bLqgFqj60QMesAskHOYsklWx9NBzNmA268EC+483htaKQDLg5tMkpr62AC
13PonFoeCqQjCjfeE8OpdLr/8pIvhFjMEx674VYXn7aBtrDYJl/r/lqV0h5r4Y9JdXKG6Os7T1YW
FGUltcnz7DYU6fQsRrURuYVgoqbaaRPnO2OkThlrC5rPT1UHz/DvnsgMhxr5GK0I1aQHV58ik/BJ
KVMnHtkN+341vtMZNufFa+SUj/FDExlbAKEoC1mv90f85ZgVIiiGl9leig37K4ALdlOeiFT2D92g
0aTWxfzcm5kJsShqR3XZpaWHe6IY94XKNWRhtCBJ+4TQe1ueuCv92uj6SJFh4LFfMB3KlGQuGVix
ZmBr9t6yK1BTZqDaFZmBoalBwJ3x9qZiUjxyEZdUk+3hMDL9BvIAK1Hv/V1AGEo+9YU/lxlKQWef
GtpZlnOKLTIVBOg/vgsd2u0yWLgOmRdSlEAbqMQn3Yu7/PF+YIQbnhIs6wwwYWirvXJ1hVkSiIDp
/X+WEDi+xMVh26KYF2uwLvV2JLrEmbhMXjT9z9Y80VUH5Em8Flxw+MlIZjzracFXz+c1zktnOM+h
lQ3dN+g9R/mFtVtltCETe+9KwKMSS3r7LLybLbuzTMBjvYBPzL27HUSSmbf51B2yH0yrr4mjwUtZ
Fg157wWHL46yOJcKDYKJmQk3h6cUh36v/ZpyQ6PYymovaT6zilIngTbfteX46q/WD3eXfBCXjTeV
Uul+bqbhMzqcY5u+HAGkepzEmui39ghO0+xqiVTeVlmV00rBNPCndL2hZSqwTqJj9jUhyMtrFhDz
fKB8vD8snMmoV0msdbP7LltOvzjnFur8GYfR50S4YdwXuekxg9xeVKjYB0qnbf9ZuuS7VKil5Rt+
WN60YrhD7y9b7uCjA954bRndsSN58nvMKvMTfCEIQ4OgcZDjFvE6WMNg8uJsIq73z7eCm1uwcI2z
hkpKrMC2vmUcSVumesqgQ0Lr91VTbrOX3/9QMGg6jgY7/ipC8Jj4MdgAKZuzCTPvhxcnvm7l9kxb
eAWp+L8B5s3l71e+1eYVJyM8tY9MFsGy/MJm+TWmwxMsydvl4duRXbWNisABzJbuHywIF42V8L3r
t90D801QAvGNg/KfWZVxoONP/cAwtanVbIi2oJ9pTyqy5ZWyGd+03I3gF61DDFwo5/kDJB+Vk80C
J8EID4P33OhiixCSU0vy/3mx8u4zjJDlCNnfGM9uT29UEuJv9UZlvoIe9SFMF2gQ/UTx8jV1+z/S
/Xtauwp4US/zbAZSe8gKx78a09zGu6iXVfJKdUhLsX5ywr4Pn4BChjmrXhX35LUhBCIr2a1BF1Ib
cKJi2z1Nq+phMp3hFSb22oEHnxDe0GdpUL46Z+Li+7FQOckMequ3+ATG0zrCSKshaWj9VW+94Du5
kf/dYQDRgjWXYiHB7HnfwqDtz4KLKiDtRZjstMC03nmW3mf5ckMbzcbJVFuuF3SDCdvajBxm3oWe
hNkv+qRhlWfju7pJXE7wxiydwh3tQ50x87vW3YE7fZrejRM7kW8JQfmDQwcUWXdZUxgXl0QKFppv
ktO4ntPPX4YO1FWKBjMuCWuuLwQ8qa2UC4A+xEa9AuK209VPt3Bfkar93U1G8pau0wfBKIf17OGQ
j6hINO0+jLVjSEIitfR0ck4OMDdjlkczoNAj1FDgKFKvY9CfJXO89YXp8B7SqACjsG5aiaoWmFO3
NYq89SZ1xg18l+3mCdqiF2gGRxT9vwWZvdvz2gIJytEBWFP57Xb7tnROhWc6uonAk2TRdCUOQndC
xwriL3FzSnLNKV1Ell9+x7iNt5LrrnO8v9gO+Nr2J1VDrYI7iXkwbEGZ+Fel1R96yvfYCpMowx7I
y1SQGrpd3wS0p7tGcGdYArxNTglEZWUurtcwWdOmeRVzRabegSwzkCzdi6LRsFVjalpymC0VrkEB
/uv2ScFqjDnWExI/ChqYfE+rBfaaYhFDGJcBoU1Ue4HgZaKaP7SDj089pZqAQFKjoR8VcUew/tA1
SzH7K651103rAm36127mO2a3TKnhrPGajd95HAenCT3IWcgo1uX6h92jlZ3lb55P7TjWoGuDcMR6
c8076Y4kFnd+W8Oy1B1OZ3As2vC8iEDqke+UcNA70opD4XSCO6BdhJrHSQ5HoG45to7Fjnvhx6Z3
E9nfDTI+MIOwjOaXg+3mAcLAqydSAkvGK7435jfs3TfFr2LXlP1FPN0Pcw3o1crnqdFapHPgxp79
wmV7rAaEHjnP18HPkDnCht0ux0uSXjdUitIU7ie5GtO9o/PFJlYVEfxi3BkxXvBOxBsntUlx255F
/GJA4X/U7LsvyQIbNVR87qVXQb0on2F6sukHisiQVAfEZLN9qmBVZSzk6MH9rtcwwhyYbEk8BCGJ
O+FV0UDm9OKMGTiDlZCg0NOcxviKz9RTDQVM2FUrG4T5IsXknMRR20N+vVncm56ZCkEcqzgor71q
ARfn9nv6aQRHHD2b7ZOccN5lDEv9TCa/2RzdkzegcTJZZwkAS7jpt4haaffjNP4j1av9p+ByjaHN
8vw6amx7LwMA4G7pPZjdLsCMZ5QHhZ3TLCsfVb+8LFmdNJrNLhtDsUWhiiHPb9c1BBLIplpqMSbq
9dlgKPMgTZCsGUEV04jyJYLPOYi1dgoYjHmiyAUFU5HfCYLs+nfMEhXa7VRuPKXpg1GIbquot1vx
M8ilFRxcYL2JRRFDdDXGvziKfpI9D6PhZ3Zf8Qc9qe9+rBd1zeWR0u4hKzkIVzpZWHa7wm12rYNc
LKbFXKdBqBHXjYKEYT4oN35rlMyGcXwEI3l7MRBSdYK17fKGFFJioRYNSljZdeWp5TRHLQBLSkDu
yI3YrBgZFH64tB9OtTgs8F4cehC3t3L2S3S6WJhPH9S2AiFmpF3YdI0mkH79vVypiy4vbFjETTZw
Pnpdr7DtdOztY3+XfC5rdUmzIxBZefAV2V4OkPq5wrq7wkON8WZCJSq5zALF0T35EdWy00SUdoXy
DQovNHzyJ0up3M+1vj6i58p+CeEYRmF6GOqvV4xc5mFlt8Js4k+oICiFqvyBHKL8OAmU60J5/0AG
QfGIUvjHMJJSYqjWCTUrqoOKaRG9XYcZNEsKd7Ekscm3lE3hU0jJR/GUx+Dv/t1ErBwQe0Tuklka
85vOoUsYXz4bNk//Vt/HMV/nl8L9h21sr14R7qKll1W3QZpSxaHxTCLxYc2u3hAMjBMS9NcWa/ML
TsKetH/QCANgwnlJ+ABrC7pp9t+hCq+Lz1qVW5foFHpngq+ZccAi/8/c0BCqrNGXiSC6dHRGE/TS
0k8HuPVsKsUN381LDgarIgmJD14j4U5ZnRak3bDNTNuTSNZLMFwrEMxnD0yryewNB92Sh+qGSwiO
nfprgmEmQMCAxTSCHNZ93s97RQrjqKGxcUgvYxeGJfTn5Ag/rNGjNUVi7ch56RV4CNx2+c3+oZVo
8CUkIcCrTRtFVPZA0/MiSXXibAcsvasShvnKBFOXhMd1JRiulwDbIhnk3f766VtgYs2zag5oJzcJ
tj5T8URSGRL5uA9+yRGCoN/cJfAVTvUTtDB1wK1JoVzNxo7hlABN9HjS5skuTW2n35QUBdnGlPuT
pZnBEsep9JLE4/QF/uCLjmuOIhx5+LqeJQnIW77AgY1hY27I5KP8HwiShUPtQSRkGKsZygi7JLqL
bwY3h5vJ2Q/7JhlE2TR+W001HbGCicQ4qgU4uc83hesobOl4qNXv+0GsCE+QhWpUDBn3DwyIhv4H
K6jpeDmFMyUHettabFdyFqwdP93xA39Bj3UCo7ULKJEPmKahKylrLFu/WkvKrIHA9M3RrRI6BaUB
ilChADcizRoQe/+z5spth01EU4cfU6GX2rb2876b0ZmLUgU9A5Eqwz7HKkVTf0XrGgNqXtCbFfiq
53N5LOay1TApjnXz1X05M4W9b/jyKEgeHi31vpR3MGPULNjZN1j5ews7zFsIJkNiLlfmU+55Ww3e
aiKtVXcrU3mqm9J7m/+prDEF/20wC+5TMolUv4gmVfBXkKi9mrsri4F6T6EYKoCIBm5k00/fuDuh
QcGSqS/trmj7g0hxnetiGI8vbdapBiSKxLVExQNMwK3qB/BNWBDVnEuarQ4fQubDJjaFqrxu3b7B
ywWuYQvWtK+XSMQtCqFdTZsf0iWLb3+oPpFrDjY3G/rlDZK0i/7bIPdnq1NBbhHxYjc4LUnA9O69
RmdAY5fxACbSjZe021/7satfTsNzW82RZssYnke1VwAA6CZ6Da12Z7Mt0J1bxu2rXJ1SHEqVncld
ztb29WSVAurzQfyoqNIwr/Y91cvnYsHwQhm6CLhOtM4Q85nZFguwa0K6Tv2LWQ68Ev3oQnfGWAAk
LSE7BIEAOCQtHQKOfhffR++dDQwI1N+yu2SfnzgssW2k3YtUtpH3GODbJsgmp2O0lSHogHLh/LEp
vn79X8H1wOgIddSQLYQFI/zkHuY5p2zrJLxPlYKOaItHkRfuVxd0+XygL4TNvQhMvrMpBFJADTx5
WUy8bEF1kWR5mft+RXEQcf08lRb4r9MzDRdDDPVAu9RGom/PyxsmdVsqELssrAEUg44a2JJm83ru
5wsfL8Z8C8iOwdF37G3ViBpZmsHEjsCA3ply/XU71YBIRsUVO1OBI0MivhrGwX9q72y9zqL+MvMK
swpMdDJrODCQkoiiEQ80B3AAMBRu8qR4dgDt1MJu+4lJR5KCD2Ie8JzdYeQY6f4qDDXfSMRVDek9
uznqBGEvHjpKjXn99i/AN4WpCrzd1FIbztu/zJ3VaLSP8+q2SWVEmVVsb1UE2XWvCHF6QSrnC06y
24UWsryPqUQpLr5z4fDu7BVbgoQ38fxul7y8u0rcSJE3HAQD8mNN3aZl0wNtNRnOJ4EiDvThujGb
6JI6mfPN8nCtSSB6B4vI1YPG4h/LWay6BONBJ4JSP8pL2THghe1Kg8TX1sfawl74rfp5wPbSheHG
IGIAAVdH7E/KFo12bWEbrA3pdXUuX752qnLJckYhR9DH3Vr6NtSgF0KTiVCwD6OtHPBOlG8sQWPn
q4TNWLDr+OvZ7IGwl2ghgIEpeMokEw+kiidVv+rkkRbAZY+swbFDts3VNeh4oSptfFR2lPVMVMSK
DFwKonGXU3xwVp/60JNQqRxU1pMiXcjRso34K+hz++X3qkMl2GqTx+wUAXw3v+rIVzBo1mYWrDPW
EfF48PJZNh6gkv7ijZd0NV5I81FoeW166gFReHd1cLgcxFuVXFT+BtEKKLPaDFmQKx+wNjkEhUhY
PHJSpU9krZrvMaYihJvOCFBqXdYFNgyfDZU3EogbWvs2++xZBeYXM/JxIEIVQz+F0np8TCJOLXTM
50lugKVSVJicESiGiCZHc/OJlXsk9ZSOQn/y/RUmNTz12Rcwr0y71g0N404tXYBldxmzfMGsSK6W
aWTjiLAOUbKUHjflibDJ06fkZtwXzp8UbTmI9GmKfACiCtGYkLHeqXUpZmuFlATUecmGAXk9wZj5
GKDHk2Y55u0cbBx5Vr5WzzATqoJFaR4Pg7SNszF8eBcGWq/wEF/eUpd+QBIetPVMbJ+uaJ0+wd7X
C4+fCztidu+Q5lvbCkhnnJdUDlOWlczF/eoD7lN7ucTppRt0LPMTXXx0VICB0OrY1cMVxsF9A4CT
UeaPWyTi7N5oJ4dwCHdY4JtNgv4eIku3e+O6OXkBlLEZabSl7VrNckXhNCOLDDNEM4FnotJH+e8r
aVoH/AAWSkCAY4jaCFyEQihTzwZIhbZJ1XP8FpD3VncUhKaf8MeVOGPDl9chwEOwTiImj4CvXt61
ofOitdN2d97qK9PIMdZDtshmALb5muwqKYQQygfVucvwQb+NmdWUbc9erDHqS4msH2gAkPNednK5
yWJTeHNZNtDqBEOXnEbLjdmsymovMeI3DzUXpcmIweW03PiGM4AShwzW4Npx6KQfdNZlQO9Gsl0e
fQ3hKLaBamc3jebAsJE5Rj3JKg6J4ubjkNAjCddlqVCdf+S/4sSt38k8WInsDteR5+Quwu4znIX/
YW5VO08OoM1Y1w56lg5eh33f+vp7nvbhy/b3mkLSzMhEkropEG/DQM3aCdl7pvIdeDbK0YqsBGwf
wMm3QHACD+GbEcncGYsgPnuUOPzPNz9adJygxtgDOtJVGrxYvnIEMRddzQlRUVxZVuo17hf4xi2E
Im0uIVP3gQkIILr0F0zHRT01RVHuLMh7TXHA7w6sAXJQnUgBrReKCDRtgqEgbX0+uXR+VCKNi8ka
gIWkbscPcQKNAUaCg2dsoxPUAm77HJi7s5sQk2dQKZWA3BRKH388C7zcVf3RX1EDGCTu/zRmuNc9
q42kQH2FuN/uF//el3Mger//quwfB5f0acK4/LvlQjMy7lA3m/8CFYtBuG2bZzgpDJhn/yIgNX2d
QillJs8Ap6FxElN8Zc+qAknMdkxJInNVow8S32Hya7QPlGcsqD5succ5paLZvMCVsYDelc5c+UJL
Z83gZ0el2zr6ojboLqQ2JHu/d3Z7H3wnc11/u+IJAHKTozx9kbVvWuTiP5Qx+eQ8HihZRataZzGc
u0KbgzCepJ1dUKfGjnizZSfeMQskZDbBF7pyRRSy6JgiLHMSRXf5RxhKKwI1L4Tlpij3LMouHp55
PYdEGeKmDK0bHHZYJcOz4Qe7lGbnqSf9yyC/8kMS/lShQ2ePB1arfjqtLcnv6+ZanHpAZoK2IwKW
36Ws3Eyg7uRPdIC9WjHoIcMuELKy3jrjHlI2Waioq2dT+iOPxYSE65SR/3K7A8fe07BIe+miYibG
ywkuQa9z23Tp1sLJFjM0srYnIz2ZnsaxMscPpsTawRxES9ypxOtESUKp5eOvOOAsx2msgP2KfMWE
psYrWzqS2CN0odkrnlsigiSADntx5bkRFr19mO9kss9rD0RfNZ9yVf6fp2bg4zTI5GxteKdpOpM4
+o1MgDs0R/qZ1gthGr7xTR0n2UCyJrYkWuYuOQtWqGisqiQRpmgUQ2rJJ05aPsNFvwH/sBwWcrY4
8EKvtMu7qspbNm+K2rTOrVBunV134iwQt4ETMOBeU7NiaqjLp2EKXXpBPHuverhLfGPcj1YshK/S
Ug==
`protect end_protected
