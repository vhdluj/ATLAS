`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RtEhbuHKmh3vAN2BFWN7ITXzA5h0499Z1Wxvu2NX+gMIQvrK2DASnCuzMbgNK/kQuUDvTzaeG34u
OtD3bLJMKg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IzErDl7bCGIisDvOSbICGQ/PXdBQWrvxLpOIEx75Md+pqAPBOQPpbosvUGFJLy3XmkJgFH9kPwJM
+bbIg1L6JkoNPjKb2xku/8VVxenG9wxlIns/ZvcUPFZ+En+Awpr2HH6T2ydUMOu+qjsHh4xb3v/x
JMuGB6nuU7HK/qdDHaM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ngN5kvI95wn0bL5RoMgcdU7QoAjRXywJD5bYE4xgjtFREszSgQ1yZ8/iV6H6OZaEMyS05TuPG1xS
hFurCNao28wBPanjs7TqcyfVMw5Uh5Jt6Fpkj/K4OTA9SqP/wIz+1t2T0VNpMZtSNESIsQai2dkW
dAak03pYMtgyckKMbfRBHDsUGXSYylk8bsD5iXn6A7GhmCPs1EmXs3zpyL97xPEFocyXlditalOT
oMqfau9d7bwk3icL7lvM5aKMcX8WHI2HUUpK8FoSN5JhudItss3OHzAcPlDa81y57ZsgKiOKhgAZ
4lGUDUxclb+KGyU9nkOh0v7+rr00V5U8axCXkg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nxRk6jVQEgFbxsZcEhUyOWgA922S6HJSgp9Q1U/85kAdSgsbkT9r8Og2qEaIS827H6P8xAz4w2+g
7WWGZDiiNtc8hGncbnxg4sqUBo+exieQMFG3KG3SGi3qJXnnWgVIykH4FWZ8eo9P+0ikJI8Neh7X
TnEbBulwT4IZgLFB9mY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qegTzleqcxC5msHpyfkT6VLmrbHCWdJQtKeOIIW3+B/cGiVXBvOdO2n1gg/SXG8qPtNfv2hff5JU
ie/2LM7pWcDMl7pwmuqd6QdD4wzFvcnPOoeDwzvgCqmXHaUCLtnBLKY2GhMP0N5F8M53yUQflylI
GvNM4xcNCKYkNaAUjyevXhJNjiBF2tnJLcmkey1+5k6noJ7kkRRmWKXJY5MFuLYt7ktiPx53Xtb1
Txi+gA/ShiXyloEGhSwKc71hsFEn08omR6Jmr5q4TDDho38HNPWcoq59CjGddy6gHrXD/KucckQ7
hbsFnm8r7PkAAY+qgrJy+LjxSQb2tjEKViApug==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28400)
`protect data_block
DmFvlAG242sROgooVIEwiuYqQQjwkcylnCJeHrMrnRXmBLEEUrScqO1yMRtppBnwqbI+8dmY8HlA
EpXhLb0m6S7X3CP3lDAaj8UHpf5N1iFLHYMG3j2bhTc/CmEFGUeyPu2gcoNW46ZTmrWHR5TqaFhL
RxwHmKuverPp5SlFOW+phOJvlGTetHiBENj7W3ZAAw2jLY+SpmNo28L75zDctYW9bMN5mhmb3W8G
UOvZS+rubVcbT4NxcCmkHgIKcK39HF922XY2cmdufG5Ena/Jn28+/lNqidndn4ySZey7voD8MCla
wrglfgh6tEOiZTSkgiS1AZkpsdKLGg1aD1lzTgXDCuP9u1r64vs26tyIQDZ1b+C/4EvKoTxTxhcF
G8LnJft+18EeB82oUiFk49+SngK1cUUDl68VPurNXxI+XyWe++Hi5TM8jip87Hk7au6H5N8/v7AA
e+qk2dIe2HldMcCigs4QZ+hMf0Amr916RV9wdN61BkcAvbzG8oTNeSZgHWWxlZOrJpZCZoQ8oE5g
Osx3cIrt7Or4MJYooMhgUYAUITFywZVu5UCe2Xi1SJfuipuSzuPKcpV5RgjX2rgBeaNXb0kpUkgN
6nX+lhKcZeRRItORB4CuATjaB/DMZd9KVyLDBJhiJ7Lre4enKMJfBifHMDX9z7K2CuyValbOzYAD
5dvmfyeli4OwpEoJqEW5ObuU0GyEy+ViIUMckvJ5ou/yb54Py2Tk/EI4iEfeGzz9l9pb729gBOGo
WfjWCplhGMJTeMAO3MnS1D2g8R/eDCxeRIy98QoDKMhZ76lQgTTCVdZZSKLcU7KsATtNhdYZ62GJ
3gip7GL0u6lZjsUeomUHqnAoeSm7PZu0Fg0b7RGLRrDaRgRfLIYickaLeytOaGKzSb60bx39BGQR
iD2Z2zmzueQmInvphGi2Y64AIGrZ92qbx1jRv6LdydkmiLYIj6Bg2gyHBpi4Qxj08lpG9ZwIyYh2
h7AS6cCGnVzswz2pB/ND6yHSHGo/E67RY9kWzqltIEYf2ejVVfij7WRd5Wmpzjt1Y8CSccpp9c/O
saSNGOaaOglSfIWXwqr/l8ZKRzl86X9WWI2oktYDZoy9v2PHge8mnhOOgBo5JS78w8Pe5AaDs0mt
bdhU3MZzCTzTXgNvpS9Dr1LQDyBdfKDdBu/r+uBchPiIRZ+O1zc4Lz12hjErV456Ij8J4Indy1RG
El6TReypNK/G6WqQ/9BJG9M69+31+u8BmK5NIPC5WyWZI1GZeETomntg3xIP5t1KdMYdvOhT6QWK
jz3qR+vPnoxLAPKEekkqQODpOqr+GV5SGD6cptTKKEkJeJBM9b1KuP/sitXiYTXN9du7Uw6hkBV8
Jxkd3H2fjFPnYg3LwoNloIt9lr6dw5eCMXirmTKNtLa7DfQsAaV9llboA6QQyhFfcU5ywQ0nlkcd
Qfm2Yed85cLIOAtjmAeXIPuPoMp7HXWVB0jDSpII959rmIpKwlv49jjHDoIsIGe80H1P1+FjNx3h
NaU/selD9ZuAYQIqyKlj43abMM7QMNMFFeyXBuDx/y0ZQWDnaby9BszuZluHiLCiMil77U71s4Nf
oU8CaLvFDuyAspyQwLlpkZOGhKQKO5cNnYirACyeTipJ2n9thSpRgBMa5/Cn89rUENj8oG7rpODm
XxNg4bxv3HkfEUQjbBJU52Pf2pF26t71Mj8DD8xdQkd5705XULM96Ki2K4tnvmbZivyLE383B0B2
MoJgKaj8FTYHOjRcHJempxjumgT2RofylIbPxqk1dSdKQxSRsKfKlwD2CRbnj0ONLPJvlhfVUw7N
i30tmvtHcfSjae+r4yx0N99hNuOVlVYw8xYZGRVs4XKr43R4Wq9StvKzWjfPypVM4kDr85onC+mK
dJN+JuzCM5KL7sORs5DHKeJjtG4XNwWbgiOlPZq6FcOgRjj2o9TE8aPiUfEU8f830tZydQRzedzF
pr8/L509l06eqVCpID8SP2/UVM1CAj+nieez1IP7j9i2KCv8/D75R4+lRA+6ELsz15ZiO5Y+MPHA
jbumVZf0B54fJGCGt1XPh6SWyu+mWOv9pnDvyLTeTd7vH8Dc/FBVNrqH6dnMIYRLvJQE6OQcCMBn
Is0ehjuOehfV4I+LO/BUWdejISonwzLP8S6hqAvayFcllf1p58EOYL3OQ5aL6D9Ed53wcwWwQ5Iy
JjMqeRF4pyLUB8F79XitkrEyrgtm/ezf6G2wBlNdmynoNz/lQvNBiA++zgjNXRyOTAYqI0tfe1GK
otswJOPHupBIcLJf8p3GebaPrNJdhepgJPgSj7WtZzyTZN1Zo2V0ujFQ8X1FOFAa2psgqy2TA3TD
z/h4/x89u+poeF0lRJnDTlnaETIJW/RoFMBl9IXrfcbxZwjDqUtY5UUUpAlbT14hLq0lugEMDjHg
Jl+D5D7sp+SghmNX00jPmlUYFyC+5bkRRFZJVQFelRoKe4YuGSlwjAPXX1NuKsn2Uf7so2Uy4qEN
tFjXfkett2BB6t+5kIZowB4zdufEZi3dGipnQCsQ3edm2Q835aQaGvjTZXGW6YlrcBAUEuxeVCnm
fKBK+/iT79WcVRgM4TnuaMx/69t4sFtS3y0vW5O7lYEo/XicwwcHUONZbLWxR9UoqrXdJ84bJNdx
6eispSo+lEr8IjLNP4mkxsJk26UzpE5VbkMxdzHu/uFvwLLOINuGBq2RLSu6qkXQM1lbcNn76+NZ
ktvUKRTrLJGQcIMphr0yK77qF0KK9Us9nCrsVptKmFSwjdFLiZ/q0fxTX0vfcbMkS+oCubg0PpF0
B059LwKJ2h5bEhIXhVbg41GgOk8g3XM4dqcBlkejjufIxfswLDNuKbQwujlH06bKWfTiNzotBADx
nF8ONzXWc7n87Jc5F9eorQsHgasP7VwqCZKgIs+1xYH2vgr28qMwJOGE3gRTPG3+WlYRZlxM1+il
FgpYhd/qhS1MspN1U0fL+DrHTf7qYwcMoZ1inKzR3a1gcGN+1FETcYCxz09GhcCnoCLzakUymE39
DMmKlFyKvsJ0GNGZXOeMlwMdVo3qmvu4PRxnargBnWhO9X70k34AVIixx1ZzywUTJMncw+HtuivL
w+ZilDnP3WZEeeVYGP1QA/PVU4+ia7/Vz6ebm9g0R8gUpxdlp+GnCqcyNq3G/zdYLlJYAm5HWfld
1sARZKkcSUiZskjWbWuW9DaFiddRCVVPGjgjkfzWZ3PV2f8m+RxP40YsbgjTkUbVzRkwejX23B0T
OPcITCYohi6KOrjFR6m3B2howptmjnmQRVeXL2TyfXolcklxSnP2g4sIi5Xz/xP9nKQKi3ed4J6g
VuhldwN5UTd4X5eyb2AwP2AzrFPLsPqZROwajYSZBhuEMcEvlfRP5b0IANOcwGz6s7wNTfn8118O
gPoXyuGIXop2QUqFmVf0RH9ua+XMI6HBlhMZbtcqBw/PACeOSFmBiNTpmJan6Yl4KLyQhonCQ6Pc
h+JUsc1q+7aP2e84a7TaKMU1pcJRTULEhhmbCwP6pczBxrpjRSK8zka7WDrl1VENsroGU4jS4Qem
G7jC/rW7EsibkuX/Zex7SGvl4SCOVzlqS69VCs+ZRTJ8xQLj8eZTZwlPjHMSqJaLb/mVdkRVCcY+
5YXT0ag4GcyhFJ/2+hd8VYM3nHsjjOReOAloNI2u9bzVwr922loYGuhLh83aU1zmsPIa9OW7x5hr
YHQg98MOQBRhKM8zmJc9q0lZSaPSoEwlgBMgKcApJCP0fvIWbHpZyB2sYx3H5Zp96TjpV6It/PLQ
lNVMvH0T263J6PXwVOs6Va8Ox4KzguZByz6tAx/hCCH2kwdtLzOKZdke2/O/Zp8SmQFl6F06lD6e
2wowRsqrSUNOVgiBoG3iF6ML/Hrz4mX2tBrSCeVWRnNkZZGp1VjH51w9svJaiqX2lxh95PEjrLSC
fl0MNzAignU+ud9hp17L12ldPY1VwMDIvjfMD+KTKzzRGthdldF7AROTFJwfgBboO3PGa5eEVHFi
cmEUaUWBJ2iNeLIFxdGTUDRNpn68zU7Au2C9F1WjSoRCV3jXnMW1O9oOZT11ALU7jl4/uNr/uIUi
euCjyZKjrNZk9mroyybZ2VuUhU6BNCSTWvS90hJS4NTOEn2/0vbgVbuU3BPAYxp2o/4AiPN9/H2V
LuAhSGCC4aWpf3vKnjiYoaLAE7wTAgwmthEmArPJoc0VB1FbAzE3nusf392SlvjnwsAfR68XUnaJ
mzj64e2O4igry/7chLKJJYvEsoMgLo+j8nTKtt15Sn/XdX8DyfBkyI53tMvqS9I7eG3ypoz6Vhau
ATAXAZG1W3dDHQ+qjSa742sCKyMSjkytQ0ESAfwNWk07Yi1q1AKUKO8hHWEuon36kb3p2PDJs+pR
qku1YyNNuMh+Zf07qEFktYOo1pRqC3V09e0mkWXoANXtsypilvP2fxxO9NEKt8HvkqqU/+HRgOSY
1LT9J11PyQXZ/kXOVdj8n+DtKMV3KxGzFzB4E7jslRAqxFLqUznb4kjmiFn+QwK7kbUCZaOuKOn1
uP24HCoYWfYcGDuGeiiRN66OCVzxmObJ1J2hZFLbdcoR+6tQqcEqtwnYoHUQOGhqMfvHTm1RqS9/
n8CytisFHs5ekSdJMPKTUpGjDThwLJrV+4IBnK6OHb/AS4mbD8f2EeIs/zhR52tt6FVB6xyvwmU1
oVk9znCTIBGWbv77daZGSWLXdvT9P1Qyni8XVtayoC4WKp/bNgGeE6pD2fH4a8PdB8eHBPq5nzgS
jWiAaL9POS5GkqnwDGlV8KEXumY0+tCTRb6uHZdxXZBiPCr4m6P4gaBvlrdm+kw22s/SXHRl2S2A
EvWrlOxz43z0Xs8X/7ZxvlpxjchNeCX80Uf7tAXzh8yCgpCXhknzaiL+JxoWpseJ85nlX+vT/4Yl
hIlSK0mUNlxfOlSE0i6kvdjSkGhdv272o1hXwSwDvWHaO/rihgIv/qFeu6SwRHWwkx6G6krPsUQK
Z7l5bZ/5EsGmGHupnt44EjUyUusdqtmCae21Hhja985+4u4LvIFe8xvbYZmZU/9JwJ4v9tajmtqB
cMhhoCAvX7D4Xw/6fPfX51bQkoLubyyxAxtPEC7BfxZSKYXFqSk1r/P58h6ghkK9sFUKMbwmkwjo
FYCR13wSs81rBrDLqoBfLOoQ1mA9jPpo1O+QlzplMbjnd+XTTmP1SHWVj8G/i5iFxwg+BiKDRRqn
N7cKo2Ov/BqXM1Yq+yGQgGsfL8gLEXtidsUWr19kcm29P16sf3LzERrS1T724zsLc+ToPKTmZEDh
yag8YRCAsGraOENrmBXbeE0CTDReLm8hNaD3sYby0zODI99wg5yPCEhQ9ftfgih3y5Sq2sBVY9sO
QAxU6fjRM4KhpfTf77PhaBOI5tAzdvIbH7aCU6z37b0GjCG/53y7YKW1xY+f6PV7ACsbkonOaobE
VcqGnfLHVlCLcl9A/nFhp+p3LGQ1bQD18cjjuNAsN048tuoXu8dA1cNfKM7kAuVEOBae38qs/g2/
e3L9KoFHW9yt6o2gwdE8/QAGL13FltyEhIQM8+EAXtlyyMAfva6HSbPyksxFMQWJzcDb0TTdOqZ3
pxmlwZDxClIBrJ7sMKt2AOxQOOQ7AyVp+QsNOYhc4kp8RPv2jl0dupWIz9NVwNnkQaR3OOtquJSH
0+TUr3DLvnFSMoo0uQT/p6r6Pu1eHWaSxd9UUlLo7irOmvXxUEfuJTghty6oRlpZ5IjT7kIUPxr/
AX6ReAqhy20+ZgP/Y6RpRNcXFUAeESDQvRDLZtPFWzLZvagSil2kIzdrDBv1+XdO5+E8xr2bMt3/
YpxuP/tNaMwT1DMQYM1V46C3kEdXsFiy1mtJLy7jFWpxNLul3gkTC6hy0lHucNL3VZiNWVvIIBK8
2dCPso6tlYW+0vVscOGIhVtPgDr1cEDY6oGNN7tUDWasfKNyL6PgWY6pcRT1+MIHPiQk3ozww0hd
3OaSJQWaBKqLmhnIDdtVMpSBSr4PpuG4s+ZZn984wbdItlMw20+J9mapYjLoW82Wrf+BjSoVp6Ib
m3923C0qVF+8XJb0xvPsKHc7usVy8GYKlMg/6Cjbsj3JJjky8VTqZDBq0of9HbIUGqgHT6G1zGWC
KzFMSss+ugUO+ZFb90xYdqV2rncTmj6pzFBRhlA9PKHGXZgKyDQP9CwRTM/jrpqVwXYx372ilQ5Q
F+XGJbOkqDVNhDf3bv80x0Jzw9hc/Bp+dDkE6e2Vxagyl1te70+KH6Z2n986BctVs3RXwab4WUWh
ISTNG4zj9IGW4q7/LGH1JRfMJ/+OvtW4ouN0E9HQshzylvyj8tuM4NVwoOnAFO6ySfpuSo0MflZb
5megZ/siSfAbn2pPBecIRWC/+gM8WCEjfwhd+hTN9HinZlu/8Bhs+5YPzkvfmEebgb/aab0w6kH2
eMsiZNrm/HGTQm9FIOJqQZdYJ+Mm44W+HQXI03nS/jOS/5BW5k0qTEAAX6egRwwLs/1W2jOc5+4E
WWIDMkyuVF06M8Qa4ZySM0jYEJdzGfstcCAeCuZ2rIvyZgrkfCQm3k74+95KsQnCj9A2QmFWK5In
afTSPx4j1fyXEHJqBwy1S8Q3FDu0rj3D+PIAsC+YKKgRAMcE4pCbSEee13tte1BqYBiuMr8AHQXK
b9E/BHGRCffLJwP8FVAR9iYT/gwUShrwfgnIBKaYaUI/lRjEOvEm31yh2BWMIn1QldLPMEyViZeV
WGb0AIGLjM/Bli8FvyHYSI6g0pPv3QfSo1EYoz0yK4ce2yCy5cX79BRRUtk1jnAQCCWIoYL4bTT/
O2Ioa6EZ8TkjAAlxfwI3Tu7I+dBNKLEsSiRtUdUESoM7lel18p2yO62PahMStThStWUzyn9rDm0m
mPFs+VpTAM3Ra3Fo73lic06Nklu79EOGFsIJkCqnUOgBFW+jrF4jZZG92Nvjof2ZA2zGz06O6aTm
KwCbWg6obqrBk+rl8NQIgEzf2JbO8RdXeYaqR07WxnEFvbzHNMBU+2SJK3VsgG9EioccIwI4qi1o
t0fQnS9JExGTMmrC+oYN5VGp15EvicqXSFRcOWBB9Oootf0GUaRyqdHbShRG0hXmxd9cOVXFbfYx
ibKSJIBATKY3QUpfVh0A7hYBnIy7COmkhQ1vIXcN9ADHmYJBh7nQQ6G1SHkn0CUnVuI8T3x3jm+a
k2Vy3FgHmrQDYGw988CogmnpGWR5tk5kYbvwhev3uNj2X/Nd4seusKGmgiNKxEVerI9FId966Xr0
h+3zT+fSImtJT9HBZd0GKAoR1K/V3TyZROGqPQOz61KNEsLvfhEE6GXIovh5EuKgM0QxFZMIbz4w
tr4uvbyw6nvAZGKd4k0Ykhpfn2MoTQzP9o6xmGvQ83K5O5nM3QtBka/8hclw5Gw+UPZcDx8V+VaA
9WAh+lE9XDNrqNCQQjO3lFJ1CAfHd5VvqMLR/YGr9Bs1bJWNjmMsM4hVeOOyfQ3UgeEfXkqBdFgR
7WBqNkoBWIRJZuzyuZr0wm/dzIGC4Afu2OocHX22mwBvzqbjAgoOp0q/C/ikZ17YSOCmnSAN/xnZ
OvPGgG1gbwir7Iu5RvydLV2xrmUg+VnWebeD3Om0xAGrckQ3Wbkpcm0kCXNmDFIlP3KVOxEFlbBg
AxNm79pt93PyAv0h6BIH59g/BNICaTCYwYMvQXU1OpxMG0hAmS9JDvF2TxruPwu7JsnH+X1taBTX
UEjYaE93HJnqUByDyvZnWoHHXkBsHdn8bsOHYetCjcLyUulinFND0wdTf89uFeoviD/ClYIMMJ/t
QR4Elhn3uYC+/1Il1ITr2Teenr47ZACLd8XDmR9QkTnP02ok0VX7Lrog+mRuIJJFHjPTGQgVZPH4
1Eu2azPNHRkN38Uo+raJTombFSHsWDAAVq31fHwxoO2bMrmjp9dWbstjHalWGJuSOhJ1yH3M/uXt
YzTcc/O14wsvfeGNzhza5JIklzQMcmCUHpdhjIbhHphIKYlEhGxULz9hefFMGL7C3drfo/+VP3Gx
A3WNDKh7Wr7v1AmyTZpVXLzF+T+xZqIQXHlmMMNP/jUJLp9ZuJuTskj6vmcT5fZ3CYJxClfoCXMt
3M0EbEnfufqdLBd+7oTh9JZOB58l2+cyoJVzefGA66aYjoSN0o8MFHEGyZOUyp2zAVVxFHYDtzrl
iP/zYe4H0aUQqefR9NM/odG6EDonXCLvre0eyvG7SJNFTQuA49tO6BmJBMyeez07DRnWapIfRKVZ
X1gBaVhWl6FMBAkPMwtrc5rptPHEFyZXxvCM5mPIk1HfdwgSK0QeryaeDsjJQC5OyvBnawx2xv5A
ZQkJUORm49e0P0BLgi/MQoFC8fQzZq43VC90cWLhu5x9P/DofG6RI+JuBb+KLTz0wis/bOnF2MS0
n6g3N9Ou98hSM4v/llBm/0c6N3VBHgoF7hRoPuK2pQFSie39+VwIE4xR8YjfH8kcgB+HV3b8miL3
OOcLp0apsyUmJhj9RQ0HCoBVM5zDYIiX7ZWwo14tGfGsVzmG9lr1sDhC3itxhXmML2ENQ5/JLTnO
MMPvdaySmvMSmazhnYrBd5t65agtwgQ5ewCKo7DBTsi/ncedk4KpnppFUfoBMxEQYRDeVdvMqQsx
6zD1FlK+moH9UUPWrBDa6yWHW+Ap/DdARZ9199H5yG3DQ0Q177ooFe/t6pWWsZvXLL8hAgbkf7ed
McQ4xwEjo+3DqiTzgPyjXN9cu0pQhruGaq9w4wPCeZahtlzyLy0xXIH6dO08QzMEyV5VBy3RSQUh
KYck2EgSw/kncdy+LifbhCXbZtXdPZVHbadPuzeoRDZvhZjplpZW0W9eHCW3r3PJuvFmYCAT6fSF
dp9i6Znz9EheKm8RXpwqzUQXL+zFbByG9YJhhm11/JW4+KL3qR6p9Yi9dArnyKsazJfFNLYbstid
80cydEFoTP8YpSc+d20ZIix2OS8Lt5mU5I+bzNsNpxVVVtnRV8qPFvIPK0H4wWHZ0sEHMHLsoLEe
yEl+91EC3dhwqUHOLM1ilW60IaUPDl05h6mGu3aVcx3pRRiEbHUW4nWA6mKtRg1Y2NihND/uhHhZ
XwQPyxxHdYuODwdwhpqSchaNmkAnekd97zuignWYnVnl6zIdwlKKpyCHXOYYXqIbZeF1b0pX+qB8
uV1WEEJoJGX0iewg56wI7zjmobNDNIpgmwfUfLuHIfsURvwHkHzph1auBkGo9h8KWK42BnzDjUUY
luBmsY/qJkFJ2zdWhG3MUlCAgTygTzNDBfKQ6+TCkf6sqryAbQYSUiwsL+TZYrNpfdnlYzZ+o3Mh
dxcWSpf4EIWg79sp79/oYIFP0hwqDYB8rOXamlsFfqr8dsVn/oTqIL2haEkeRYkKkLtT/ri21Yg1
od/Rw1E1msyo0IRo9+9QvkUnZvRXV/c4Kl0DODRp4wgUMFeVAKRVqZP5jEQeI7g8ABpsPPu++2P+
0TBMXJNwZbY2DK5pudLo2If+5zAzGO3wx+hYkpRpaPtWloe6wApMVb3RKmPzPMspFy2z9vC0lkBO
0obtcXG6kl1278hnVVQo6/d1jYT4x+x3/vqCvH94QVvDUe/yckbn2vJh79fO1vY/03eW8gFhKB/r
SW075g5atkDpfUTOFjsi7OWbjNtlz2q6X8YGFMHuPppSJ7fVK4SH1tzL4yF8TtZ+S7c0tEnFOTDs
3gdGi5TZKDEZQzKH/NsHkrUiwC/B7rMMtqaseNs7UUq4J2BZK/N1bo7P5hyA/22lQqbiT70/xfDO
i650P59QxZHf9CyuVsVYVGJoPpPRpBy3AdkKMtzEYE6MNoi+E6waAsmFGkftAqlxfTVddW4L8JX1
TyjRbN/FjxUVS/q+PIJGClELC8vI90dq12hnTc73+EGsEIJw0kS6miAUdRjXIOGsgwDDbee7F6J9
R4Bv5jBmvoe6eDMYNkI9sN9+M+6OtWvzKYfYasOObYSxpw2CccEpKdlVB0m/3wEDWCyxU0N9zClP
qBHO1HiQ154PeLB5seJNLDCx8FICQZK9fdof0necXAqG1yyA03Oz5DsH280od7oKfqANGgoqwpMU
O/ltA49VMZmaJYRXxL3F09lwteSmOngkdlZfEIe9bIZhu2tDT5jXLfsIOJMJVZ6JiK37JQpzvKci
jkssemO4hUPe97caQEb19PuWpWIC4zBaCKXwF8954ee/D/+Mx0In44Yh6bjYcng5//rcxEv2G3zN
JmwiafMm+1ueF75Myh6976PoxHFA9rxwy4wG2tL6KIHubMLDwjCQRHV2DogVEBWWj8Qx9iRXWmqz
IsnQOwgSYDRxiMgf7dLnIRAR9fCRS01Z1+U2LGx9Epb+lDD+nNwYN95k7h1WiL/ifdqX1n+GYtXu
9m74wDjBPsWDerGIBI0EqZNYmn7zlkVLjAL8pfYN0duIRFHkPsUrt2u2wIrp6XZqPgk7DbDTZyi7
m9I5Izyo6L6EPxDDqBES+cDVCeDt54QmRw/yn6rChhOJoO4o+SH1uv9RoItc5G1YCP72FsWF5fT8
dhOS7+lVpzZuxqtBq7raa7w2GisGfByNd9h04e++TYc+fXp56Q75wIIRtNw8IuyYtH1Tw1Wvb4j6
d0bZ+WixUcdNntwLyCqorH1axp101JUsLo05piMJi9OZ0XzFIgZDJwHT4kXjlsgfzjwkZcGksidV
ekemG+VNvU/TAbrjdoomtMISo0zUT5em9AGjhkrLv2gunaZa19vhiJcT3khInZR/poi+8CmQKeGF
3IY9mUTwKm7cYm3UezSFcTSknYLVCiSpN6TEPzvHnF/SG5LTswdbhMlHtFl+VPziI9GoBYxjPlUE
nELc2iBBdceuzQ05O/27blr14IugG/SMTLa0vUAIBhCtqKOXCpmSzUEZAj6QcHt75UdPiMV2T/ZM
e1+lAZB5Gc6ZhSaKIHBcBXTZtQhrqPSphuIUU3J+D7onsiu+T1xsBRcOgMtzcYXa6iWD6C1IcShk
Gqcp4lpvFPxq5UH+ThWymsipdn9Gkhsr7qCjfeNVMr/0ZeOMPd04Ojw+z06s3xLT1PEjVm3ERZG6
1PNnFAQBQwjw6ofEiHtnqGAROqz3v4CUOXpShQuCf9xpYqnCjoAGhKwrLDGIIt6j1qMfNQiNGJsG
k/HTAAAgZwnaWkqTzNuvuxePb2Svyi+gBdLlHy70Tmy8h0aV+rCfNClaLjrcqzGG2+PXA43ah2m6
DecwCHBUok1fmGweJ5INDicBMPO4dxWfKBSgEmHA+7yIpE9NV09BbtIe7LBKu36Vzhjv+Kj3LVxy
YNfBiZzuFLhH2Kdh7Tar4x4naNU0yJlPHcIU8x8h7fDIE/0Ooi4OBPA3hMmbp/u9Wx8x3GLQYxHM
UV+XQ4N1FB7jPAVBAZ6MQICGv0tHAAKfgqo7aRsAQe2w9hHjjV1xx0wj9CN/AXyCQwUoqFAe3Ieq
pRTyCWgSGVHFevfn8zMqVx71u3rV7kBOsrgpTOsYKsGKefpld9hVJq9y763LMn4WFFArSOa0IeE9
d9zu047GpLYrJV6efLyWY4DCHq5BGZF5GNbA1CBNtN0/2rkrNoEwFV3d+rh7ZUgc46MxdZ82beXU
D8wDCFZrI61ARZbKoLkgCvgmFfoPnpQ0VwYlmU1FPFCm/SA3S1LmtrOE+lc5FRcDNWFxXloyHQRJ
F3XpoehDKegwDytRhFwelcy5MXGPjYYxS/XaY0VfUnxOcUy8oM/k6L42yEXxN2lPT77vtHpzRHvg
xQviVw74o5Zx5BDqsky9zBwYOrcJ5x/l4eP165I7m2YGQbmC0v168/4BsLVsEc96hLZXwT2Gplp7
N/pi6GNoCYFeUYVhJflM8l3WLitE36hg4Bbr7yzrbmE/BZa7+keuLNKW0Stf8qJelAqyotZGHpnu
5GdXEP+Kko6HQxIikz7NlRl+Zh/jEjfyTPLFcDXo+YAQC//RWF+z0RjlkwSk9Ax31MYeVi4aUWzW
dkZ/OE7jkbExRqBqKDO1HO+oVoDYH3Des3JTnenZnET3QFzPpjf7yYSEB8p+cB/4zjomRX4yIof/
CF6YfxLkSVaSPpsBwAln1dLUqXhxQIz2WIlSmlzoW8hMQ9nRUOARRxrdIAKQyaLeO72NY783AMyc
MhYBcLp7azgkY42cninnQirfPsyMU6ZBWhKM860GFQQApT4ltWaeAyUTZo/NZEl7KFzG1ZdYJDTN
oKzzjhum1WoZAMYU5gadSU2KPD6UcHBN1mQnIEJ+agqmP0xoD9Tjio3JJHr+qwTJoQBaFmgSD3q0
uOa5PH1o6g6M9caIgDBpqjsjxFZauOEXkdz6+DcBtu4YRXa8wI3VIJvTQcGC0yRqM8NmaYLy69Bu
h94QD6pFLkeWW4AT4WdVWUuEhPV405z35s4kMOfVcqQIHjcr3NS4zoo3h7Q/ieiuz2u1QBH94XjV
9EJQGsw3qB0CmjBDo33wZeEIFY4DsYaqCYSh3Tg/u+pa427hlObQV2WzTqCiiueZs0/WQKWuM07M
EBPuN2IIsG3O0mTfIT5KHv7BVZObhtWu7cYCwjs/QrtMviOM3D6AJwTVaXxKXfcvLzxp/xQy4VyS
3++VBqwLiu8kWl8GoOZeNPLuoIlucZo1DIQPv7CdKcSEjTi9RPqfPYSgocgPq76w3jjH3shKE0lP
plI3/JdzRGXTp0hmHRciftlaBUG2etScKV6068tGhXjkkHsbp8d56sITbbdPXoEn+iHPmG1tYI/5
QmpuxiDyrvcCEZaetB1BZSRgtybzD9kcCwmJEuiauPOcBfuFnFp5Fktp8//EPtbCzwAI0Hmd4mxJ
AFL5TxUal2T/KvCA3CovSQ4KoDUytYtv8uAdL3mQy1A0IsKvNjwULhqwMx8nZtW+oW9hol5Q4JGS
EC85qp9sLnD5AGZAcDF+B9yp2Lzn8llTXOE3VPhQQ7Im1EypwtI79osV2XVG77q4AU2xqg9LnOzQ
+sGqaToIwk0MnJ8DhOFw7mxIpp6VKW+AEtsJOuAPbIwGSfZLJ0DlUP9zvmkLu7FKD97KTWIKI4im
zykutrc8fLMExVm6KBvPrAjNXIsZDNTitD7UWUJ+jZI8qKXW6m+utk0QzuNv6nAyrw9Co9Pn0IDk
C17XWQ1ikgsZacoA6J+reyE1LcatgiI8znds/0Qzx1Ezji2wEMgMzfq1VgE69HamyMF9CuU4WG5V
Pe6ky5hD4RSAYNVfvcogORJRIuDIgCbBHATmog9Iw27VgiB0sJJjyZjJiCzjSVxIvo8Gaz/saPkr
An+SGNCopR3IZhx1phePaPDuwC5RXhgdZPRLqtiig4ImHoSR7OetORlFKA376UCahD4tm8paBXp7
rjvMx9HB439rIKEIc+W9cHpARrQ6+Q5ZhMNDeKRwCXtXrkFbXK+OI3c/w1DSsA1qzaIzbWhdOece
1sovMCS3qEvTVKk6/D9jHFBkphrW0bvXZEPCzkh68y01ABptWaDT6vorfwjNBga0/kkPNZwG3Hsk
fUgeBkTbb5t8ICr+8kssbC2N03JFVJTd0UHk05nGw+8GAU9XMczAmnD+h8plMLgHzgpHgZSyHKy4
FwhSo4sfg5/XoDM9fneiz7+BjpWx9uLggdGV1EPkVXbePcvI0hB9hARMZX4LFJKOoylP7fdSPmcE
1pXPttx6C6RMwmq9LXeOXvNfdIuwS0383rVUD1Nc0QvE2j8+Xp2ITTcONGDKOV80GCSf/GiVcUKN
jKP6VY8sAlKGSJL+aQElNLli5sqeHETQUXOgdSf6Mq+DZMSDgxg8E39jQW4rkWPgE/MvQejPYUkp
8ksQTYmksJN/xcs4cad71h2UtykLN6/C4I6MxGsxmX4sB651uYluFJoYcDBF2lw7ckWRamNY8zAe
Xii6Spb/b0ZmY5+ipq6277HP7YEc6UoxaMAxim1pivOaxfgIPNOZX/1H4C7WPe2QIu9bHNBbilWA
xOHBeBHIc0/bkCMd///xUO8S507zU3bkZsj3oABbzfHYoM9LCInrAvjbwPnD8PVCgZVONGAuCbWK
xNbQ1LtADQC9wstECBUoixhRqJqMiZ4wSYSwFtaJYS9SK/SKsamKV8+GqgGEqCdwR2QrdtEMzRhK
DZOESH9lUlqWQZt7h2XNMYtx+aFLkbS6UFZ2ltLsz2eXLNnNz9GEnWJ+SVUTNZ2am0e62plj8Dpt
auqCvLmzOA8Gi8reolSKYjQmPjrNZgKvqTLmUCb1ShyCLgmrcfmSUSUw1ZHkxL14mNZ75BEzR+vu
yj27hUzvKf85QccWJb9dyXd7BfN88YS5zkaxFQDGLjlQtsvxmDQpw6fchaSULx7HsfXpHnIEOPCT
1SuUhhUKn2JuJ4MIZrioWr97JacK4zBCfd9RlLYwDy5inlpJBW4YUdq1/l59SisPnBF9ml77LiJc
To7KbkjvV+PgNDlcCTBbV36qrfeXxCS+ByJ0gU9cDQhNJqbRsG3JpSMfjDHPdxGVQrPm8/CAXzmT
D2d3x96M2yGMa7CzCcvMFwDFl1D005jblKiYCM7qTge/WLL9jxyP6gvrgqtA644CucySLcvluSq0
14zp0JelXMLZwASZsZgkQvlP8b6IOh4vHDkV0WXo2pmoNoA97b78JwD+r96Y+Qh5QfPHFXkN2BTC
nXn1mDupbXb8kIaBXYobg4TSR3q1reYa+827nEBuFK1pxUla6e+XFYN73SfgxLF3e0J2cHogSjyC
I7f3IAJZTLkTtsWeMANni06o1bFOrQpnYb/oKzvLH8xadW5XvqQkOtKg/fD7F8pNtnAqCZ6kXLjb
JpvmG+dCdgSYQvoFzwGCQp9d5ythnIsxUohehWz+VghBapaZoCLbuYgjMCsaaPkXT6Wv0ivphsbL
tNA8IhWLZZK+Kt7igGHOhvos6aSquhEbW7iCR5V0HW2GsfFvizn0AXjfNfKtWJNUGoQBooygMyaX
ev2fpwjFeP3yb0dRLjWKGZjgX0TBjohlGQ6linCoOCBux9XctGwFVS08X3hi4kZqHafC/B3JpqPT
bSFyyr/w3B5oSAQOjW2H6soU84S8snyAvCBcr0NTK01WzEGS64/zVM1+oqzjAcaTwXOgNOD5cK+b
w/Mf7+/n0NZ8/KC09/s6ZULnRCfSRYsnFrj39j/F8ulcIj9OsnpM2kC08zBB3D6WXbag259t0w+U
F4kxLIA0NDNLz3kyqGqHmNCCS36fNkkulDp/bMl0Zmir4IJCckPq0rGHdFMjakV+NyeeZQMGFWky
o3lDYc0HgpkVr8uqT4Zr9PcdqMNg/8BxhSaFFA9ZtfLo2EWsa6tMAaXpEfFglBm8JOn9FyRf2aUn
6USEvTxTyD/WEzm1ffyW9iZEwDPua0CY8+gG5ZPokiID4UunyFX86XRENEmahNS9QSZjP4P6+s6P
qCcEJ3wa2TM+6YSqViAS5tXni5CkW0MUpXq1WqQzGmGAnjS5wWRLzK3GIa9fxSFIJRWBLgwz4BE1
UvAC/JVLdtVOy6hBH3fidziOd2NAOmIWh8aebIYJbv6banIMn/TyZL1k0Y4VtwsvaPptOOS/78De
XqKFqJ1fG0BaewzVk3oQLE+M/BYElT3RoXZ/ZmlMcR1GAvzUtyA6Cag++naKM+rDkjUT8YDxfg+5
TxuKyFwgoRQ/Wd2HCYgsIzz6VutnYC2ZpnfE+kdJAZO+98qtAAGOKPn1bim0whQ79kGDZ7haEeM+
NxNBK6aOnlJ3d0iRXhikeoJUfeAlBTdrgtYPOTBDG+8XjDpO9mhCoumjxAOP6yqtsBNbHWNbvach
4snuJtc+FiqW6ApA8qHkAMcMlFlaSCCQqMFsrOklXKyeCEGSvrQNJJ1L0WV2EIdsye+k6MppAX4A
c+JAugZyVfsVPbn6r80FBO72Vm7WCDRZXfsImczhC8CRsSmefVQmY+tXXTHRtfavdoagpE+42vhv
lu4SzgdNh+Yd9nCGf33ZkZX2fwcJSqgXALjRlpmVHNA/U5wxIl7Imr3EJuDZd0bwGxSEr77aZWuy
zKbfpWnYXlXbjYkGon9n5/nF/vWk2EwIOqVCkhiCsGwhn2wE4U5289rv08sZEMqtHqzQcoKK+9u2
Ggg9suulAjHD2I/1l28SlAb+sXrrvqSdZOwwXBMQBtEaYB2tyrZpu5ZTm3QUMj/5CKHcN2b/BzyS
YI4CkzWS+GvwQ/icY2TVf1fgFUdwz9LWfmQiPEcxVs4DGjvS+u5CKl7U24rpBEFiKSbY44wEdkW/
SDdZxQN6WQ+yCcEhLgdQyCreL2cSgUIrxs1rEKBtDUU/z4/YCYWSzeCmKaBcd09it4STHAnGfdjE
XCN4fyIAJi9rkICMS13AtCYCknW5K1xVXmGSSLHISAmUpXmu8gNFLBOk7M/aNITSPMR14RUHsQGc
ORvycAXC9NLzclDLLp5L4vP+nF4PEaUO+4VegKTiaofnOU50K/8dXRKvgTnh9B9U3gpTHXqMK269
h1nDzhTpX947D4FhSDazFGQSjkKqovsTG+yHTcARZizRWdLwdDXztNoXN0WPpfNK5soJyLOIdSal
/3zT5Dd3npKmf8zRxCWVBDnMUNVi/LGLo84J0NCgS3xd+bIBxQ5iA5qHJGXqSV3jNnfd38vqUbt1
LHceJPOrB1cgtNbAt68W5Y36wI+wU59HF084tJQOTFTMgF1Lp3OCTSZda/0dgnYyGrN2tt0qVFtc
yY9EjnAsG8T6BgvLdTpnejuxi0OrP6zG1HH6EP1pDZZz/liNFh+7ex3/qjJv6YnvTbFk2d+IhVU5
IQBRyXA0Fc624B2C7KR3ae2aF6d+treu16qyvQmhEBhn6ZI2H70Md2IkLT8svHNlBJmnVX8XM9Rd
uHJ6FC3vH3VZ7hvyYXyFgDj5ZrJGE9+/kXrHxMIwTPgFpiZulXbP8EOC7B6ecKZ7c15pyKDDt7f6
1O4yfwaPW8P+5XMH5TG4E+/6O2o3a4e15t1wB6PfC7D73rRcy5/U/pBi2d1JPAFODiCoQamJy05S
viEbVifIySLBw+CFRshbN2g/e8x8o6PPHOZDxWTJjGnHLf+5a5R0Q+rRGf2kn6R5mCTt1q3huDto
S95rs9V61KgeuHPOmBHqR+yJeN9Uzq4WJZ6qXEZSjE3jP+iBKkdIcmImApeo5KQWSKYi2LtGPxJx
9N5X+6uxkuXC3TvYoRiwNbRqhJ+9zmR5RjVwqf/cyUXVwyYWB/5S9xGoVx7zmlBYvutd3wOTvp0U
H2EnMI1UHHkFn9I5lUIzx7/OeIf0bVuMQiCgtFyKdTEmw9pnMBhlZYP3itUjEE83yhf1Ppyb9pGa
dDv+fPUeRbjzjc+lr2w5FX524S5WcCAOMqBgObmc3qI6/zTstVdLULJChTRc7KZ1eOry72IZ8ou5
x71uUkJSOefXIBrK5SapqNZr72SO0lH0wD8L+icZP38fRd07ZgLFxHI1Rcd26Hd99ZX865/Gv3YY
2AJkwKHOuOBb3XNHD4vYNmkjO2n6A8KrJCkbEopuwQnXODc5m9q50tnf0WYBriKk3neFaANdg6ww
/L7ECuYf4D3XdV7mWFp4JH7UjlnOXh86UeSmWY/dBCILVO+5ix0/3biVFv2ukydysE3G4XIaPef1
Nzt7AxmKnEqW6D5rY2Oz0Ghf7hIK4O19Tj6I7BU78JPv1cark7kXGuY5pDLO1IE4r9ZwkNrA5ROd
rE+RSwobmztXBKaJYSkmQp41Vg9j+5z41Q8IWsui0D0CoXZLOvJUfWT4GI5kxs2cSh13YVjx1tV0
stJkkji8E43TtwvgWgU0d3OojmWwT913kD0PAQbl7oBwIb0uHo0ozyZujJmmYxIB0JJhtdbOrNjx
KEp4IDynbP3tTboNpyZgSW50aqoQU4axxasgKNJC4dXi0av3+ksKYyCE0p8dqEwnFQX4NuWlDKof
DmOGdHyh5piGtz6kVwMkXXEBz8xePO3zXTAN8/TyKvokgwmm88BRF8WBkiff+9SIxiDpX83+wPnO
DHypPdgZLsq7WoORn0gmU2MB+nzzW/v5fqo7dIAA/n/uE0SGZt1bY4Xk9MuTtoagRH4HIsY+Aqmk
yrpwSdMfmIasGSCYG4kqKwqmaEacoHl2gmgoUDrYIbHDNdCyjvOeYfaz9hcic7xR8jlJu8l4wq3X
1FUK7fsW0E+XlYlMhZC2IEe/bnUri0yUEz7F5ovyeG3cUdbJF8g6Al+bKDke0MdFyTGdHCDa2Fef
Z5MCLmmtLqMY3xfNB+XIdUgBeCi3YssK0rpw8eSU5y1dg4ArLTF9zufmtbo4aUqdvEyCGuhBF0cX
7eh3tpLTyyr4O3eFKHRsk4krXwdcRdbMcw+tvL9BtR6Fu1BjFbjVCGDKl8ohi7KUCeS+s/B2aY00
w91LxoMj+AgGgWebjISGxaxvflFhsMEXUerEkaeaLsL80yeWXOo1R/C1gS1gBJQ1uiMfWOzJ36oC
L9VaNVibpurbwYNnxuD2LfnMkXJOdiU76IhxEnfVg6i1ujtr9kdoZ3yKC4DMPYGyJY+CJCYBh91K
DHVBYMOoJ6PpAspxdQZdqumEfCA4lGDSAzBeHWPvn1fOBz8rNvPvjyd1eMhjEilArXn6NwJGfwTt
jnpg0N1ryOFzwWPfORLJhVQivdAgVYgjVRz4syaG7w5AopglS6DoYLJ4lRtNXn6rRCND6hcm9TrT
gQaooO7gCvecI2vcO56MJADMD5CljP9T+I/xAlOg88u+OjEikevWRTwzs4fWHGM9Lxju6/MmW+24
fonwPenZvbqP7vegEIgahRQ5o/kIRAukv3BI5DZxxAAppGcE57Q1moeLKPPuG1RViB8fXiZd31ow
B5CEIMuHt6hxsWUuUy/i2i9mQ4w5s6pn/wR0lmQVanbivOuTQ1HuxLPQZLS4plz91A0m/5yT3HAn
XyceJag5oUKN7LholVsYWHs045yQn1jgKnXfEeSW0st5DZ3+g7NaX+yRbjpm8bRzfRogHWOL68Mu
spp4oEYhOY5tQ/e8WPqkwnF9UR/b7khPOjTyBQi0eJQ2DkQ/av9jhWIy8w14H3WT8MsT47b2MP/+
5/G0MN0vDHRoa1ApAaf4UfkVBIkOYp6IVL7TM5QISGDSCQK3KS3KohDnZMQCwbInghPbGQgoxFdX
DmmBLDmqqbQ+LEK2GDEYztyOXzdbjQn+vp0rBBOyc+MekKKlsB5oAJwBGxLywdCHkZoC4zUZ8n0m
p7OeLB08f2xhXTCNZttZ6EJgBt/2PWE8CqyFrj8auu7XWoD/KACeLtImyDaR8ZJfdZQCaJ6OtV10
I3RlzGSnBsgUSBpMTrzI3PO8/BG0uR7zQTrBLabDoIF3LX2V6JMLslsdFhzOF6UXqPj66q6q/xWN
DjyGmD5PcM/ztH05Sg7Y1mPP3bHsx2ay7pzaA/0LsX3rdI23TVtTdtqx8VyRXxi+We3/a9Vji3HH
r2EroMTscraV9vjZHA5aWigxBAop9ACpYDmnznrIJ7cVkYa5InjRSz3LLZvSRhL+XqeQHif3S3XF
dUA7/PYjTRog1zY+EyiJNv2CETPhoU91CdXbJLAW9ZJWTXjCc1cx1ZffyUtE3E+xRzEsBo8Ucc45
IoNPojjrBqQ2z7tfdWDKjv2ytn/gYPyoeCG9YFeVrN+mQNdmXlnf7X6YrSFtqcEf+hgIy5OygSV0
jcymAI47P+SG4vhteMySyLSHpVkP/ClwDoNY+ewSmOSTCvWRKl/vwfBClcAEjKN5H5dfC29h9DBL
tnWFGelBwfO3kxqxsf3Z2xgoir6i6muO3QTsLxlqWaAox5MP8JxkHwnUw1MXyHEUDfx7M0sCwuKz
igei5ozWceB2bxtdDCsQBubdN61eGtKTDU6nikNilQulqsjD9NYMbRb6xX+60Zz/LCi+BfwUpEvu
XesC53ds9SQOEdf+9chdVbIcLktvuMWzrj5XPnG5HPtX9vVOOskkluoZXZSgdPehYPJ2tYIk9wif
5dU3xshb54CPMYfonPQQRyFSMeShq4l23szGUBzyGdYmMBZ1dI0yjWZRUW7L/FOak9ISP5AUfjKs
MgO4Ngk2NewHXRnYWeR8SgRMAYNdTmvAFGWKEiRQ3YVmeOH0LFvGDwR8aTiTw2uxS3tTWLK0P/aT
uJYPpAFH8isA0o/WlLxFhe5IpODq0MbKsXtB473MolzLEc1d5GZ/+rpEEJr0U1oVGeJw7Kd2pGlt
zSvntqGy7f4vre6ZkfuewhoTgiRSOkHQ6CEGtf5FzJHoh9SMoxxmtkYui0ern8QlDoqrZlye2/PS
fsuwyPGNyRHF+WTDh4itoysIjHQi6JqYgp9Bko19aALwipn192QGTmCBCZrP5S0sk3jF6t3KH4ks
PMP1a56aApp/eEkHS4meVu465GxJXXDKGXeMju+B853bb3OL4cun/FeBTO3NspuIzySjbdPTs/lM
WiMQmqiIKtQ4E3HmIvRyrPK7evpjTTgr8/9y9DO0C3DLfERAOrTAGxzvmGp2EufS2wJUb22x6huT
A7hzXKL2oXKYu1S0z0QOy39x3/1yJuR8wuGjGSVPHbxdJlHQs6FY+6S4CF8bJY2pC0yEZ3x4uJU2
/HP5+f3Ufb+GozL9Tas7k0rT7vkGbsBZpBQVUka7XHKxT2iBxLXMDGwiUy0V7Bd047qGEUxk5G0i
TjdvbEfP9cpwZmXajS3G9LhT9yEwUmcVO/kBlFGcSbCVIYBjG2jbKgoVhHkxr/qrHt/nyi0/EWpz
Mu5azI9i4O9zxHDlYdtke0l7+t/1Ic/GT+CHG0YhyH1IiYhctunoLVP+oW7Fy5BCgXW9uyUZ6s6m
9d+8UPygRHwP0MKE6v02PAQh0rENcP95QFNUWIyg0BqshlGRb9CKCCte5Zlcv3WYQHPmNwW2rcnx
vQchTpSb+dGpcTp5AhUe8q7dsUAngfjlgIdjqWoHDEGuSW85gfLSw4epOLHAVMOBCLuymx/nqqS7
mWyEZhrIq9BnAEesm1wAqJFwW58xedIBjTyiKqbFqvXr6gbcGckGIBLnbSCmCdNatQXIV/Jg9SNi
CdZatvxYZP/69kJZEibocSMJZwnL97Ylb+au5B3KQGXFylzTiL8J9IuyaX0A/iEC3XLXNYT1WI8i
erYqL6CuMzoThm6miEEHpAwjbcJSzcz2D3vUIQATJB3j6ZO7hmEKd9GcBMpOuJZvlQRkpIkPsA4v
3KMqqi+qkv9B63pFlHAkWtKAdGPDR5F0pa7iyvxE7tkv1/D09p5GfPgfOOopDv/L8i5ytgtPsl2n
bT/NmkeG8HFEbKA2wxuQUPduuI93ZvCryvXFAyZdYW3FmLiK/kn8m0h/HIYmHc8tkk3ZazKXAhej
6qhXxE/FOyIQb+o99dM4VtPe7Ir4NMe1/30ugFMVxlpKyhB5XTtdVsrdHubrR5+AP/wISSC2TJTc
/Nfth+6m9RCmHUN0KkCXopiHYr8aqrQa/UHXBvx94MeFvJDh5DOluZ6IB9TfE8Y6JN7QRVuhoCt9
kyS7mqpQsF2WdKE9rAYfO3SdAr2NkuJ5sTtX3F/rr/mU5kemspRbFhWsihQhL33TuMF9JJx/xajB
BHqHY0lXv2jFzHMTGsXxiDYVFQyrDtIRV885kNfCDoAnYLnDTQO+ZtsUphsI4pzKfsrLmd83smKN
FbzebY9gbpw45Zyyf+eyspgOc5Jo3nfi7IcuWddkt3NBo8SHOUPOPi4uJwOgnfO8ftyMWa6UDJBo
Dj5fqzSLfumgCjKUx37CF48g6iEJLYyZpbJiX1bDEBA+feGwjEZtdF0O3rI7xw9fQij7tel/v5mc
au4M60j5lRA+1oxag15GYrV9bTg6s4aGy5CLPUOlc0fpzWMgQCojvx+Qz6yQc8CV6fzDeXLv+ouP
ixQ1OdPjXmUm6C3K/QF6moFDPtuC3Q3AKtEJFvJDU9KjakNlyin/8MxXFOeVDcNPRrZDkuryr9SS
R2+l0c5HVePU/J+hfZqUGUrGUgGIG+/IYTqH5i0mzl5RNhGhbdFWFA+VkSHN8t+c4XITalFYz2kG
LlwpQGrRGZUoUqNFSlgh6P6V8n4T84Qm6GPNiZ4/7F7EegB3Dd80vOTLFjX6UVaG4C6cJ2017Xrj
FoNTReVY2h8hkIb2wnsNIirW7nbv3UydbSUsGChg/EyVzzKn2yPaM96YvOpGGqy6x6Cw1zPl3Ipk
c7nr1/NOxmCvugdLx0HCVG5W7gnzALXFBAyGTPSbAPvl6RpC31MIymTLc6X5MlZsuvSmkgzE/9WS
3+As+/nBAjK8H8KePWP8E4BqAt3xX7Ju7b5Z1bG3oZAVU/Rz2240KFPmp3CCrrnCITp/XwuDBXPl
RSXeDHUdy1iNjdnlnDMlwh49hZ80WNJgq2KJOMlrQLuF50MaNYnsyAq++2JztnNaY+8p5sess3wu
kx31+ILS68ENEPa/4XMY429DO0HdA2T0wOufRWfIyWxZMsi21C0pXn8sI2hOTER4xtLXCD2/X8hI
jChYRFZBFNAFNgx7gtR0P63NunG+8IQNt5uZEaWPZwzcqY73aAgl0CYJJB5R56YnTCRtKfbh2e0Y
SYYtG9Eyc5a4UVzq51ch1RO+GYm6N7JFHpnYmKhTqwpGvo4Q8UpyzWIwc89wuQUv0NMD37Cs007z
z9MRbrtxFC490o9OY2TbLkdbmMrPehdbz/hb98O97iL1o0ICalSetrlMzI748keLIHfGAkwFVTJ/
+bD+29Q0isUiX301TTIPktCvswZjMLc6XMdpLyf6mUqXT8GmcPrSg+jFQm5QJRFbx705JGzU5IzT
Fcn4Tz6a2CMoOkwhJ1r0Bdh5WuRkYZiTbIroHUnv9WxmWNehuFtTOcynH35LhU0S6uwl8MAJ1AVG
+drcGMo6PmhkW/ss3cM8B475t8o1tHJ18Sjtlo3vmOiyh5zdcCiCAMJi/J/VgtAb7b5tl/euzFNE
IF6KgkvOFMTuA28dbFZAPXs0MwaxK0BB21YA1T3SL8Qr4Dy/W5+2Y0tkb7W2x6GzUbpPXzeID4nt
cMS/MGOEd9Uj2eMmx4yEi3fWUnK20BVVDWWJeERYlanVyk+xhjdUQk0N7M5nSQ2Nr6y/eCBy++eR
wfmsxbCxT2PJK9QOEAYuFeo/t8mtXzWEHHIDHvky96C5PaU9gYhC48H9BYOdNU9MW6licb2QV3p2
CX2P9Ap72udpn7cFPvAJr8WyBKHYtmTg/4L4ZXzmXsLNPF7bMPVv0ybznsbXQQaUaClFsjR+3mIj
Edaqa6AKrru29BhPn2JIclzBLyKiYQweEDY2GKBGAeMxFf44MKRfBy0nMNmOJIupPxsv17Vy3K+N
3AbhlBdSHusu8O+R/RB+tUoD8tVrTXjfJJsCyA3EPPU6AM0sROBHdtbdxjzz6V2xcBXdqyC3mu+B
Qc5KGZBKMAlcZ66JphJG4MRsluHOIOffcWOSXVDVIhvKPH2wpAtBBttC0kXW9hOpGUBn2BbEGyRo
SEGiQ6osutErJMRu+iaI+KHZPUQxyHGbMvmPqmNP4wQjtgFVqhZ+sj7sz+G+IVrn09+iyF5unbI0
KPDq8okzWwRAS2ErWGvTAB7DiDb9WitLPcrELiYfMxYR/fpk4Uh0s8em6W/zrjJ0MKqAEl940aAv
cT+9knKlXG3i4iIqt6HqTUSztb8ketgoRFBgRPsgaY0XqaO+WGSYjh19E73mlXwKP+3W6KFpgIb/
grNwT61lEOZNRG8pdRkwWGKBGmHBvJO6gYRTzLk6jJmMvrs7mHt0LqfMmG1MUSuuXpW/OWgUuy9j
0JwwFOORDDhQ1a+vAdeZJOkM2y1Dq1SSqydWmJzh6Rhlbj38s68jiTWF5MgNL2myB4mCxtu+lpln
D99vnRJGsoXt9GZaT7iTigKmb7dofusd3+KhrdY6ToZDWwMXiuOxZEmeB5FpJIZ1gcLCUVEoOyda
zc3wJrs4mYhq66FxVIEf1yom7Ktpxvv8gTuhwkCwjSrSsEivdgeKcx6ImUTCJfqPu9/ZPi6HzD88
tsIaGuZTlmMAckKgektEGpnU4mCrVDnH5r1Tbku/EK9kvPTx4xO7nGBh6cQH/wT9G5qdW2BT2kn6
CRHNDFseJhaoji8WpFGGWFyoh1ViDyYEi7dHeixeUTlJ9pzF6cga0Hv4g1OCblSRSoKykDN1X0yB
wGfyc1XYgzJXpbTo7jyIDhyHPQq32qlA5U9Px8B+XFo3bHZtZxyfrySDDGnyW+Fm9gmkqXSgM0aG
pBxyyKpcp/mij3WiV4pWIsHOhmHoZ7fMamd3daiz2g1VCnTgsp64js8xjAVYdr+dHTxz8xFCTA6z
KK61FC5YWE1xQDXgbxFgUMZ2A82y2DL+LcEOHXDgjgBU4pP4dDc3W6RCoZQ+CUceyRUwj+ro33HX
qMxWJ11XOQVDCup9rG4tfgiSYtw0UiXH3aF7O6w9mZT5ZYbFpQymu3v7E2HH69uW0mX+iwXPDSop
AbJzNfjHMKjrTuBlek4dPo+v1mOJdiztax+LWrXs6NVCz4QbqP2iG9GiBhwtF9cNeAl1H8VZq/uT
IbGktcpZmj8CTjCcDTIDyYb3LtQ8AUkhAjlXoL7/cf+XMRcVUhgoXuougySaaS/YQIsVqhXKhixk
cUAOxK/XgPjy8SObGgPK61ayuScSEX1tBdt3epkdImyxDyBaUMH/Cbh5I6G09ZhzVXLLowg0DdkW
Kuzr4sgzhTzCqfg2QAlKchtyLnFUpfEoo3JweOJ9UPqXL8wnZe96+uECP+FR/lbbwSMHuJQJZP6v
w/aOv2CQIWTewLmo/E608xxxnmYRag8hYyRjacFMEQHp0E3hw/lrHkTXZhAqbE5yWW0M4Sd4X8hW
px61V1yZm/fKdM44d5zxhpR8pbmC/7efUD6B38cHbaNi2AsaltExjNRZFxzKtGM7tiR3XVJZA26J
0Mig1OaLcLKeeASQeOKHW4umtd8inrdoxSuGWUffC+EQNQ35lu0p7HGPVdMmGB3C7a/RsssEGmlO
e+FNSW/aRB1p3brNOd6sF03Ln+BiBVH8IGdyU1dMMx4jVsZ1AtciyuqbVs2GqTJ1jyG9X2cwMgFP
aIRMVI7xsT9j85EtxTOSL/WZujnjj/QB7DIr4mNFIBU7+HOGNq0lvM9/fLbs2+huIjKfhxHA1SoG
+MBuFX5e8w70hrglb6OCavQmedzoTPHhBoS9Zs+0WRzVnRSA5b/JKnqmpzVFn41ZUD1ZXZYOkoo0
eGret6Zhh5fNBhGPiAinSdeDqf2vyjHwpPKf6iJYuANIzurxE/Fd35htEOkPwpGcp+MbNIorb03D
sbsHPYawSYXoY1QySDo9rKGMfwL6tEJ/t7chUX7C4l2H5koc2zwh/1ZJigh7vKOYftkg2ikE1b63
lwa8qXSfzj3GKCwD0S8gANmfNcxrh2rs2xlrUIpPnJ0ac1QO7ImbQRUsetAr+0EDFPFQkZ+dfUhc
tBymGPfCxJMEDhwu6tmeaotCPvtjFxsxjSsUAOd8DC3JVDh8bGcIh7NvCE4vX3iN/zrTTWjByNn6
DQkX0ApGK1+zdWNyFO9HE5OjISNokJ/+PzvSIiX/uwx0DpJPOcqeenSneS0UYCXlnmeouKnMQ+I4
8dRW1j9G39yvhbjJRNd9i9f1HV+xS3m3omvcNjzmdV9kTNbWkOz5RM7tDz+FT567iKa2fTRwBiN4
UhhuGFA3tg2OR8q36Mhr2ZcKy8etiguA8us+IyHaYWnGYWvzTJOxm2oNqexI15nN1/ljULs4nhyI
j75YltZZO2RrhxTKAmJsLaua0ejsldLovZeHXNRAuDzgeDmLQyIXxMmA2YsRVZZUQYD16ELE3cHU
IPIIQL2jhcR8Q4x5dp8jbvwdMqsgwYm++B3LwTT0L/qnHd9knH7+VldibEkNKXWMxfjTHLHsj8H9
foy9qpQqUVVBBJs0VjmWuEH8m0hoMa2Q4OBifqoSQoZnBVozLUke3sNyQq1ys2lv4GOHWT8qjMDU
WSS9Vn9gyXLY5M5B8v4PxcUytUsax/iPcLhQ6Ecd9swvXC801ipwEKqwY2o1GEZ03nWC72CNMse7
zmACDmBTLRtzSnduwfgdTf8l20QI01sm78fmZQ4nypovkMCc2pfZejQ/eXzd2CyHwNqIva2sZCmk
XjQ5vKxJGLuF/pSyYxIYDewbfy82y5dhK6b2liwpd/v2e50jwYeBE0qKIsFyHHSKCLT7wRXZett8
q3xBHBdoTNqSHQWRwmZlaS8SW7aXgCWR4PA+CIMO6RWMorfHw3UXAWnx+9VbQLkcJGlkn1Rr0rj0
40yHTzT8e5x1jjvgI98T3Mq4kfO5Xs/oIeMNCeZZWF7SQ3AappABEh7eTyU/Nao+vqgBokxCLLd3
u70chRxnnTqGyviX95M7BE7Tp9TKLuSISOOBek3K96FRG8gkBbTmDL2fEKU8Op282I96CpN93G6v
jAvINwaM4gdJDe0j2jB0wyiFFaCqdD5nzn5SP7VXZOpgwFBx4OWe14vQiwILKqQZuDjJFX+Sr7Ye
kwffwGf1v+SAa8uaIacbpBRRM23nE3Gm7fUm5bUAjnyqio/vBynzYQapJuH/J4yEI+0Vf2BCA6ss
fT1MPwOXmHgUTlKGdI4H4eBoeprHNmZBHNgG2nm8qjNyc7Q57op17yDigKtLC6Gag0bWVCoGCsBz
jDB2XUJ5ANkme5MznMDRuEI1HkVSGswauVoF1534x2xHJipthyegX7IxkUdQ4P8jQJzKn7sROguO
5BbHMm0NPhIUDv6FnxzgMOS2NqYPeGvtC+bVDV3K9+fusDEX2Xz4O3NvWqW8xZx+O4v6BzluucBQ
O3ufcUZMIf6gjoCEIXIvPvLfsaiHeeRtTeNyQkgP0oSiEMsxH+3vOkA4z20s9Aej4R/L7UH8g4io
cZNx1+XWfRyK30tJtybkT6ZoXwi5mqJ7rJlfUlKrqBDZSKV3mQeJsaR5v8DQPH1C9/cUv+dWAJJp
+1YxJxORhvaUUvmPfICrx82oqHLU2HoAWtbzgwPYvo58pjuMB8wMwh0XT+xqJs6yPxFHQzvq7rds
oayGT3/UMRJTSDUouCC9ppgBaeyjXiSG74ETIQ/VxPhb5k+Y94jmMmG8AiTUNn8wCLbx58Le28RJ
0YC6ofkI0TdISqK+nojvMwAdCq2T1+2cITvuIKRSHM1JI2v+7nqY/bWpv+7S24OuUHBLxZxWOQEJ
EPvrjpJXVvfSl4fsZrK20T8W43okjJl+ae250e5dEp+DXVtTRqgIJSt6uptffeL9ThRzEoJEgido
0XzLPIgyRuAbGbnk12ti5l1DIhG0mG1mUtwREZ7Emo65RJVU8SPzbxYzVnwKJcXW9vC7egxx9iJm
IFPqEDH3E+3fNKzru2uzMQ/N1Pu1/wati5FXqAGs0sibl0cV9mQj2Bhjh/xSLzyRrvygicHOmVfl
EU/3eHRdyexyPq4f7DR/HWYsBT8RR0HRqw9ni05DPFakxLg1biJraZixDJF1CxOXAjIxP+jl6YKi
/Xf7+K+w+CGLC2IKgd4qY+HtdU+2a76Fi+s5MKN4YE45U3YNp9j+bsjhjoW4FhVMPdagwg9BFIgg
+RUGTCSfpHOJp6ZrIPLNDWJIFS2QgGuL0uUtawOA+YuybnnwXUvZFw12egF5Ow6Xtr2eTN1fNt8E
Q/9A8nus4K+WSioF992rQ9Eh9k4Qhyk5rwmFRmut+PvuOE8oN23XieEmPp+YqSGyRlftBS7zccQh
UCXylbgxzZiuZkLgg7KVgPqsJjl3ghBMj+SjAo3t5TD/Ah069a6eaJPMVPThYiixW5kSjc7sa1ZO
y11OxfxC7U9TYAcsJy+yuo9LqhymdyP8Cfx7MwiAf9gXKVR8FFQmGT1X4ViqVe88V+c+pErspqnh
97pvA+bjYsnffgZSUs7c31l1dDdgHRf1qXmdrK/CzyZfqiXHrNAt+PTUnocxf29lz2pfU2XeXSwI
4hy+zWXTjisfi3Ar8wOuTyojHvtyezcSnzWjbq85BFNO/XZ6AZQE1CEDkcB0UQQiRUttWngjrU+u
nw9TjnN5cTnTwXKcDW3aO2fOypnd2dhPmEO9XRAkzENus6dfdgzvQRjDhqCHSXh2uU1/ejNXaSS/
SldxhIIx3CT7EzwwJbTCfabPjjYSkrIV4jRVOpRHEAmGIzMLgP7y5g5s3q+p8cCFQTbLu1cbpJ2F
ixlq4fEGsFF/2mRDGMU7YCA731aweJU13fglsMT/P6MQkJ+U3G/SU+0mrAuoSwCxb2FVD1/4usRA
VSe0Q/t+n2lvrQnPyE4Gvj4q/u5wTG5pC3xwG+OsMWHf7SbonKHYI6BHSylgQeYDM6XyPjte0xQ/
97qgF7sWh/krfp8WnMqiCriTbERf07oyAPvw0FrrVffK5CHz8w2t1SkiYFEe0Yul9NID5pCvT9Lg
Ck79PG3jrvge7ijm+AYjfwD4w1JCtACUbjuAl76iOxMjk6i9teazB6HvQX7qe6Rkgl1GBtDWPkK9
B00e0hZMJ/tM5b6FnK0vZ1N6cfAh1IwYo6K1LPeie9nHUaZQQ6oW5tqQqB7kxr+ECyPsSTEPlQ4g
s5buItwxFFKtTOdi9I9ZH4ofS0uxz5xf6+Bzk0hXJdFpoU2xStb+WDoJajD62yW4Tr8wk1MPlyNR
xs4yarHtkOpInxGkH+1OhrfyCvB+Rdi9NpGj/q0Phqqt4pTKi0cslZwNC52jk+yy1JyG+iqH2vEF
28R3UOsofFZ2bEpsIRdspnDVcHpueOLeM0kg2V0JPmYzkZviH8l86NHboec+T937PDZMS3bC+LTg
3rlDqOW338o8RtZmHVhX66YY9QC1KVuf+8ZEQ6u1QaWJt7D14DNdk2kK3a6Yzz4I3D0NMcpmkegV
JRQGVkHQLh7cGKAJqJKXodos8TEHhw/eR5GuAOYDX/81TXyLAu+aDhFqvnoL1F4MRX7/dOG+HR15
9de9fxA0/CaMbliQX6oTxh6x7hLV1PQYhUo3dhAriXIbOVnKEMyBJbg7z8YpzIgMBn4dRtUov7Ez
rjdEwkC31EOjg+QjIdkP+bsfjL0nmbDS/XksClunMJSvFsLe1+vqqZZTfhMJVlW2kuX+IDzJQpqc
ZpmcjwVtvD/XEClD+NxiiFe9XOvaU2VdNPsdQvtWWsTf8hKPWhqMTZq0RKVRx8Ki88AOh1ZRDvi8
JYEyhhlRC5rVTjM0TbYFJbN6DOYrKMakxDSplFgkPMoPTLBFfRrEbTWn5bNX/uEYfk/RZQuo9Ctg
lwr/SOjlRHVrnRsdP0Huy/HphxX4ckBhpd4briAS9PG/b/xvlnLfaLK+C9uIXbAL3ZA6cHaGtFU2
0DTkaWszV8d5WUg0KeH6j4yBt6oQ49OTAUOxkQgINmomjSw9uDJQg5tOd9Qj5dYXn23F8my/03A6
16nzDS8h/02L0oszrXRqW+GIoiij1uDq4MeMQh1DJU4WYibq+U+fS75Z9yPpGQB8AsiZkuXo25jO
/LkBAuCNr59v/DRc3rnYRGJox+uxE8GuuAQOUGBMMnPqAO4q9sQBsJd9oLZtsSn27P6ItecczyVG
rSgXUCqreNK46yOgxdtQIyxtTxC93L2BpF3dJuuGRoxnM1quCsHQfH1Vg/rqddfULb37+eyac8jd
zyUDmigNyD0E1of51Y9qJ69IXDqEdqGVxYi4BwTvqe74+JTyKXKlQ3QBsymVdP+b2t3kiJBK3iy9
J/IuoeLjAoFtqk8sfTU6W1robcBv7960iDcCY1vlawqQaBM9ZVgdqTMXn7DiVvqzaMhxJXxrOBbD
bk7Et2L8D9Rkxw4g/djj0bdJEnym1XzIkoSs7faUpWXKhVJ5ySJyNzijoEoRdUHzwPaTTfFeMRty
l2tWhLFOhUim3KddSqlxlnLaz12i42W6MIEqVmN3wDWAf2OR1+mDEfh2cutl49yP0IjDwit1d1M0
NWacI79Mraa16JXFjzOSh0lawXpRjOhSy9MhOI+VPeQUyvkJAbmoy7EiHhidXtCsF0HpvgY9U+3Y
ZruIPMc+x34syuDx+S7OeZ8uTIMMYJUrP4GijEcgJiOkZld3lIAU6lloVsTwykzDKcLAyAVrdAix
s86Msl/XOajPIagGN1rQfddfyUk0fJcqZdAd2AsLridQIjjNPpBqi4IFMs0aH5TgvuckARjVYUZE
EGg8OwbgEIgIRz0CRZShtmSl9qctYZl9VMtdVG3ZM8GwYgnhom1s2kMHi1ZjKB6rJlZrI5vhRKkd
C9QnZ0kR1v+Y+oDPQ8awoq7uOCBFclKQYtngDG3sg6thBAy5H6lUGJAp5FjvRaBYV3SWJwT4DJvG
+7pw3pgLBFki5sVVONL3mTHbimoTHsSz2zoGHj++ITlECPPYsd7FoQlVd3QGSNWGlhxSQqFStM5V
O3yLEC4GoARssIYxEd1gB4fBT4g16VXVWfztMi2ah2nzJuubNChfaLpKo03WbSSH5MN380oSGy7K
rB6k0Hesd8Z9Gsgh5F5icjcZuSezVAyGZvZ1P8WlGz8Af+xF8Q1eNOP2OeQcJNYQjolbpaWhePUe
Xjv6P4WLhAL0eemxnIGHS3F7tarLKe7kZ7+W2GbT6v0U0MJrTrzLUExK7TTMpDGAKhQ6B8I0XwvP
N6r0xZTJhjvC+18dIpzu/oASeXfgV+LYtUkGg0YGu7LyHdModsSXyHjHnq/93Zmj4DVOE+X3lclr
L6jAAgnhDHabr36l0d53BNwuEwTRO+Ui/vvxJHcOsugUx4l1EWzsokCohc9qQdx+ohpRQxpnqf0l
SGD+wwqHx8kZpBQ5QVr7TFvKI5rQ7vDpecuWgo8E6RoioJx3Km0dt/wN2yCTkcFrM/f6QI93eNbL
0gtbCzUxXHb4bhw8zQbWnB4v0e48BEVc+C013o4o8HuE4ARFe493JzUvxz342PJHQBntKnV4FYYi
Qru17+Rsgn0s78eSqc0WkwI1b1In4lVgacbJFPoKjOguFsz2sDwUkoAsijzhCdAGAljXDMoeTzZL
rxL14dvlxPlYUfecFl2XY5BQr1NzVjxrMmur8My/O0MlKaJakESEPn5QasImc6QOu+IyrhNB3BDw
KGhk4ej6QXnKs4iCcCSBxYAZ0lFEquOpLmeF27y6w/ffeBMMxddqdRXOTAjs1vFUMl8nE+8TBvos
NAA08ZDbTD+0AUe9q0AO0G8iDEy980Q22mmz/uSGBGmVinljyY/D61rC+O2xZjci9aqQKpIBoZ3g
wGtNM6C4KIi301DR4LjOZAkiU+y4mJTs9RqJA2u+zQckt+tg/orUWvfxiWgnWAN9x6OHTPbc6cDW
SWPmAvpXxcg0rpv+A1s/VI7pl/cmemERpPdJRcRWc20tOnbNN6gE2IMzA4CrxqJ5uAdRyClUg+Fw
ChNAx1Afb0ZKAZAb0WvicmAYb9uXSsePLgeu9HRDlQoEnK7wV4/CWcgqU+jN4LIezQuiraV6s6/q
CVgos29QCOuZN8h2/zA+5zjJ/CVX1CzpXfRUpTvLba6wxcUxjoYXnugeT0wrL5ylgrahLtKUqdGt
SP2C7RvJlb01BnRX6Ykg78/JihhS0CGK79oT6spNpAbzyv/QOQqNdwxxAh4tLCewlhJT6RMwirbD
AMTPh9yz75M32lvXhLKNd4Kb1Pc/rgPx7Qy7bOa/4cv68hzSJ7GZ1X6Zb0WHjK2Fg5YYdPe2fREV
j9MWg9iHe2d26v0hh1uH84c8W75ArdqRj3BDoxyYIvuBXHI4wmPvyYSudQ1CL103vzr63UhtTbeh
VSVeHrBu8BwM2fVvPViPE2LL+bjIItG426/HtUfetaXm6wigkVYLn58MtxSV8xumcHbXmDW3/Hi5
qJ5BA4Gx6Zc1xx+D8YNFl6c+IL/UNNhKpOyGaA1fciKa/UtVhzNAK1Hq5lG6FfhfoMXyN8TtQyGs
UFwS6jhzCydjiiY0dobQcMwrJaeDko0X2Cvq3jVH6nx73pvqJDNVd9N+lzZ4UmW7tinh/t3KrFzi
OBbV2uM2xejHz2VIA+0HEF0UBPUSx1V136DI0OI4pC3BvIr/GZh7jarcvmgNKwpdoQ+/XS5v+a55
6BS4X+cerHlVsDiqBS6slFd2j6M5e3hHCRXtzUhRObKueQQvCRtKyvV0R4gU5FyJ29eW06JXfHB9
Y5sQNHhUhTzWupO4ClGSj68HyFTUU4MkA7sfBZpmKAli8ii03l1Icesm4LF/D1Ym/+NlgYAEPOkd
yXiDKP2Tare65MclNL0FUtqXT9Z778PtCkLYfJS4/yjbPFXjhPRGW/S5dtOlLPmp/VU+FuYmk5GM
0GuG6hm5VmmOMXDeFD/eXPSJHapWQNFIOPv7BFLLaCDAuVTB5Ohn1xcm/k2enZUXvPgcM+LFHopg
kFsYwKBLXv3rJeQgFItIZMBGPY3riUIVw32Ac//KJ8GnQEgNtFWQdw/pVUM76VhgsCmJeIEFcVgX
d8MrrW95gubaDs44RdVjpKqfpjxlgKxf6GDR00D/mg7FK1N0rrcnc5ws5sV176a1NDAnwX9l+ImZ
XwkmeEQlXBQN14UMNtcXwSuVBvDtltrl9iC98MXornhDZARbhlimWcWUBHSdcudRl77jBmEE3wTq
p2IXNaCZiEGGJeV0nzHMq1OTU+vjyg1+zeOGF8sIW28P4F1UzvGNQmsY9UCax7BVfKU7ZdEYy59+
fydMS9d2aWSLV9pvh6Aze/hT/YhAwH/FU/yPo6mp323ASzL/89H3SvNMwn4rAkoJgzxBqLfsfGbD
EPRS4qKMzXxlHz7VJGLlvbOCSo1/l79Xrm64rrkkAtdzhAyx9BulBlvttPRoQ34z25SZ5UaQoOOU
44UxlOmmza1H27eluPr4+7THRrU0ZLyniMwycUNH8AOfA8TkH1iET92uyCHI4mbDMZylb3IOdbMP
5JtCtnqWD9Ozdqmy5krxRCpDcaEree5cejHCQEYQzic6VMdjZULxUugv4G5ct9xCNCAz9Yxk/rkN
TP080CnWI29otEI01a+OpQHS5/EwrlMRQ2virveEYdOV86yiu3H8YNmjfqeYvrw7AgMN8H6kPLYn
PeU1JvspRyL++aB2avbtz0D/ZfE2kcaRYC0X4S8VMhAA0Z5+FQhG3AtI3WsM7DpZJ90wOrgE8M7m
gbQnSR+HhMaET4J3UnIH5YKVibNJM2nfqWWWZhDilW6xCPHlw0uF+9iQptmav+n1c/5+QOAuW02m
hA2IqnD4nOpRqhb9pMxDU/eq7dIFpNMaUIWLOLr6MjoPIST2oUu74yukiiG1Mo4AnKx9WRUGkBjF
TdM9SRr8ERHCweW01E9q8uUmBdPg4JioTnrtqrwheBhb4A9A/vSNRjERjXv/r0FffwS2b8k0AI7I
r2hrZAsz/sQX1ly1htzbtt/0VQf6T72fXYC/ba7cx0bDnAHWtdyEkmJswnEqrkr5qTaDc+57LHIM
u1RjsTca6Q+yr0dP48PqleXyZTqQgRsPhE7GrtRGtMxoNEurf8WHiqQcMikZWuEV4Klb9/a7Euew
sD/Q1kDCWn9aUEpj+fwocdsftBNCCHD5/1keFddhbSqVtzwyjMqCijoCiLeUxQ0FeYy6MBvcmaZV
LE5exoKKfx7UDnYGKkq8UPsDl2wBxoBKB/IfrPSVTC46sJ6txqrNqa7RGXOk2Eb2xY2ygiiazbdy
hCbu4h5KK4F2HRiF7X9F01daDPItcQ5vj7F/RQ3hm6jGImgmalV8KpjbsDa/D/Hkh9PyP/9I6AcT
FD6nclSx/maMi1zpbWHrHE8e3czzPWOTh/vt/TtvOwnaIuzL9g9OAIdgKkpHn7tNKOzHA/J1neuD
QYR229ZsMbgBn9xVi7eOv4TTYIgmtWuKsiiapQ2XaHF9fRYJ0vybzH5LZE62gKhB3OGrNNXD/LTt
M0JyMGm3SlaSOhAlHoBH0XsmuP4fXngLoUXXGkZLcyhdJ1nVwp7H0OTAQN4w80QNWrpwVi4RyFKq
Nra6BM8dL6QjvWi3kLybygTMXv7aEZD84bkYCEru+55/J+wABXkEJTTJbBDxYCZrVrpIHKOh1Vl+
Amci5nn89kGmLLPMul/MKRzduxYPdYMKRUasB1a8nSN87y5GmYqVBwuPecWSMhaWCfxBL6Z1mP/W
Bj+8A/v4ktqFEH9tRZtha0tFXtqv/9Q58oP3M2E9BQ5AnSQVCHaGaheTM3MsvUxKNbrdduB4XF3z
mSAjHZI7im3abMMkWVmmln5tTTrTxeu0hL/VmsnyhuqTu0srccIB94ViJzWjU4fH5LGuYd/oMVB3
rxYc3gL3xv1dIfD0HfipbQicuooMyYdqzpY5Jqe7gRVI49WWmCf1do9BVqHTvWx5A+FQ5z7CGNX6
nCwtf0V/QxMgFgJBwH6CgGSCQniB8CBpaG2uUhgJFPZDr0P7+lnlQaM58xCR8tyALeJbpQZ5ARl/
hhEpGhDVvV+ec9XOuLXVu2/kxZPrFYiG9wBIdjubRznVnQs0/e6fl4h6Z2JGLoAvd9QzsvbauO4w
VvWQhqiRillFHu//dni1vCA+xfVJPOYaKLwF8fZGk1S20EqahYMVmLDEH2K4ih7VZmIP9Hl5W4gD
MO/xgVjxK3vtmnm/bxvOkCSvINCXjMRzt4Zo2Xo5JVSwZ01KuqLWT/czQLBOfc1A2BnMRvwn9S1I
3VyRfEzU+SXWtGTIURCtb2wc/N9SixC+AKdbfkbk6Q2RUbxPj2Iek3OCzFghzwgjwms0+70HOi+s
fxr9vVk3Cmtr/m67DlTt8GeLQteK4u8lOU2HgaXSFc4xWipShzN+gzv414E7zrwuVpxfayl4R5ia
F6fptt0+RY2orVEq5QhFEcAnk0ykJx97PALStp0MeZPUtW+NcFM/fTpQ9pZXL73oIP+fJzmKuR3q
mvTTjvhnj8NCJk8EdG6FGLG/+W8EozcHoET8vdBc7EE1nUGPB0F1C7nz5rDe0ayLwN/x+VMJl1uo
uyhWjVJqv1VoWL61KZ4tZc8FQepYlhHf1zeyFKd965G3zzUvkHafpmIgo1t1PoXvmps44z/6pMh4
bA7C3gA0ONadBP5fKijxKwWhyDmXvVIz15WxYG3GvQb56tH3kYiGPvocjrhtKeg5PSi9ie3SeSg/
MBytSnm36WfVdrek3hoby0/GOAzpLRjM0+v8qaNYh+RK4IZ+GsFDQWynijYXY4j0GuXbRA+7YwLc
plvDjvkZgp9w5KVlngEPrIpI4H7oRXdUWTGdT7XbFnkjd2PkBPiwThJvHw8XC6ophUrH9YWXZcVJ
iAb/Fo8ZLxhcR87xfn/XKv5fv/TZT5TiMsCSk7dHh03iIGHwI85qiKXahJCakz0ljh4xQqk1Nf5d
WPYZSp83E4AptnNmqfDQXn/aEpxum2ttL77IddwEtPIiPf839mwK73HPDOyjFW7Nbv63lradEMLw
4hBRPZug+bgEVVm5REwoPlyjbqmwfkGCzY1oZq78dMYc+AdgaUn0zF7BGWMGeCRWAOOv22sGZp+J
+hAZwp/oMs64FWC38ZFm0wd9r5/6bf0CEpmRMD0mpeg9MCp/Ck2S/46XqVpImFFauixwHT0yOdg2
8rRQDCwiFNJd8kdXrNzFrXrCfW06F9qc7FglEL8nA1DqhMtjK0eXIpmpDSgVzUXWNW0FHi6LJJfs
XHr0e2/EVLe8gM1VOj6RAdRy/ilZtBTOOcz4OMCsDEeDTqvfLHQChLxfq+a5sKSesPHzMSFE4AYK
+ezZ7uxwn2BvPzFGUBZcLdNiVbFL6GYMaXcROvicijrniYLWpTzq2IWfQlHwOLOVhyzFDrcM94mw
Unijv3fBdowqmcuNaYhPke2Y5Knjtc+fT+/0OBQvfInHc+LGOh2BIDHeU5T7RU/tg7kp9KYN0OVs
RuAUPzwrAQPvNrIQ8Tnza+kCpN/UJ+RGEoKi11N3Y0NYiK4fsnlqpVTDZEVS7JXItTj3oF8lRTpk
coOojFTPKZydIxVoamEi5R0Kw2WE/lhc3/Lwe68v+GYDMDD6Tc8dj+qZFVr1clLsaQE9hhuxn7Ez
VN1G2XtnTRKhFAFgtVAj6hUxYWta2SjMXcmp23u9XyJJVcyYWnVwYqLqUlbpGtzxVKNnK9YnxbqM
quFU9Y3znCGwLceTaVR2gC8wCAb7ElRvJE3wazPp3fHh9+fkp+K9u85Lcx/qqVQ3Kc9aEEAiaR4o
VF1iIe5AjXQ2JagXVypbJId2WAJToQafetFvH07kdgl0D6D24QfkwVOTLyVDMknkOtIAV2Unx/C6
joWfYONgZVr79w4F8KRa6WJkSrkjQI4+JeRNAM24MmKpH2wgl12nn5xqUNSET0SIkwepjOELVTUQ
fcq9RqShHbEL/Ej/3n5+jiMqAoumdD38A3nTbs8NF/5hV4iazgwCXiBKF6aEzXXZocNB3YPs103o
xn0cGLGemTN8YX5WN0+pAmPU+grTRag8JdPBMW+18lsQgMqhRnyH2bPKKxzgvdDfIbT1j+i5/Ap1
Bkr8mqY/lV0KPHNGZw0pBV8/+Dse6V+/TGMs/wXuKv/UBoP9K1EadGzjIgWugn/lmPZ1qEL7/4+F
4ERqH8tDzbGG4lFwNBvKRJH7kZOHU0gQqdp69w3XWvI+cPN51hSpi/efVN8oHgMGYbSHFWsZmt+X
bb89mS56WILOEAwmYDL5YSjjPc+9LLM7Z9Vue/SvizgMRgk7i9G6+t97BRA2AsSySzU1QzNNK42K
VtWUh6+/bCDltwUA/3QY4DURqfaRABmihm0l1QhZ9UKbDTM/XccLvzOpxtrE8Cxnq4WuOPjuv1Ub
uNEyr77orxYguk7BHfYdi/X4bHeTbUyqRx96GSTJla4dh6v3nX3uQVTZhDEhSwxSfiUnpUlSyyMW
CWdHRzJdZPdtW1KtHIsoGirE/u0mBVHfRK5lHrob5rDYOmxEOiSmElgATr1wDXdvyZj2BL0KGJV5
95xy7fZNcaKP03LWzRx+ndzEASZkDb4Ox/AWoojVOkpHHVrP6HqfUrTl0UYhcebFZeoUErOfvHEp
kkimEG0AUbeO7cuUZ6kBF9KZTmPwsNtnnmzXzZxTdPKpnuC7mICT95RDcDdn84+tl3cC2GPnbHaO
3iBaSBOQy59Pn0+uQeU7BvTqdYsLgL4W3twHjkP0lX33IdKvBwwRschChyThoBzT1b3r6bUq/Vuh
7CG1AP+uYPbIeeb+/F1VFVG3z46jy9DpIVetdzwPUj3Wj9AnklBRx5m3tBswKlx49mjn54+HDP4Y
NbAhKBu2yPEk1RO+UgH9xQvbfqI3ndY/Vhb/ZVW3tJdc5CUWNzGv4Rk5FaRdE69chIdiiwyEox9k
hySXmcnRUysCwqsTPKOdhmQJZAouhuBxNrg+fsilNnkFys2d0N2mck7GfGY5SG0o39ZnJ/l+4h2n
ml/psIrlrmXXuCHkx8mxNbqTXOpoMAzmJqfzeLyjxcJLKSeTyJlCytcu7gyJkBSYMMv/wIJYTvTb
PmRPpUSjZopuwc+U591rsjPOAizlvFUnqubqc+ymhIsYaMKfMHMV5b2rKznxzuWg2fH4ovEYNLjs
RLXOE2ldtZyHvn8IQqMzX395rCTsGpKeAzeoSOixRZQU8TCACFe0H/xcxAAwRdKZkGMjLr2wqVp1
sarGuFPClEKu1mQixIGrPIkP2PfoAM16RT61lgAHTH45GK2nbGR8NOb5GQjW8Xb4DzuGdl5IdgSc
dL4SwvHMu2ssbWVFMhDFDcfiHnzVpw334n7++rdvsuIC5PxCQ6hmgaBP+Sx1NjMnKBF34HoW6MNk
/NHg13a7+ZZuu24FOksHM+gB/8zCf99s05gBLZMOW3Fkx9GinFtud1GihLLvFhL3T6ARF/+O34OZ
PraUE2LJ/0k3LQeNH5Y=
`protect end_protected
