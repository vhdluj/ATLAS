--////////////////////////////////////////////////////////////////////////////////
--//   ____  ____ 
--//  /   /\/   / 
--// /___/  \  /    Vendor: Xilinx 
--// \   \   \/     Version : 2.7
--//  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--//  /   /         Filename :gtx_minipond_k7_adapt_top_dfe.vhd
--// /___/   /\     
--// \   \  /  \ 
--//  \___\/\___\ 
--//
--//
--  Description :     This module performs TX reset and initialization.
--                     
--
--
-- Module gtx_minipond_k7_adapt_top_dfe
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


--*****************************************************************************

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.NUMERIC_STD.ALL;

library unisim;
use unisim.vcomponents.all;

entity gtx_minipond_k7_ADAPT_TOP_DFE is
 generic (
	AGC_TIMER : integer range 0 to 4095:= 150
 );
 port (
	EN                   :  in  STD_LOGIC;
	CTLE3_COMP_EN        :  in  STD_LOGIC;
	GTRXRESET            :  in  STD_LOGIC;
	RXPMARESET           :  in  STD_LOGIC;
	RXDFELPMRESET        :  in  STD_LOGIC;
	DCLK                 :  in  STD_LOGIC;
	DO                   :  in  STD_LOGIC_VECTOR(15 downto 0); 
	DRDY                 :  in  STD_LOGIC;
	DADDR                :  out STD_LOGIC_VECTOR(8 downto 0); 
	DI                   :  out STD_LOGIC_VECTOR(15 downto 0); 
	DEN                  :  out STD_LOGIC;
	DWE                  :  out STD_LOGIC;
	RXMONITOR            :  in  STD_LOGIC_VECTOR(6 downto 0); 
	RXMONITORSEL         :  out STD_LOGIC_VECTOR(1 downto 0);
	AGCHOLD              :  out STD_LOGIC;
	KLHOLD               :  out STD_LOGIC;
	KHHOLD               :  out STD_LOGIC;
	DONE                 :  out STD_LOGIC;
	DEBUG                :  out STD_LOGIC_VECTOR(53 downto 0) 
 );
end gtx_minipond_k7_ADAPT_TOP_DFE;

architecture Behavioral of gtx_minipond_k7_ADAPT_TOP_DFE is

component gtx_minipond_k7_adapt_starter
generic(
	WAIT_CYC :integer range 0 to 16 := 10
);
port (
RST       	            :  in  STD_LOGIC;  
CLK       	            :  in  STD_LOGIC; 
DO 	                  :  in  STD_LOGIC_VECTOR(15 downto 0);  
DRDY      	            :  in  STD_LOGIC;  
DADDR	                  :  out STD_LOGIC_VECTOR(8 downto 0);  
DEN       	            :  out STD_LOGIC;  
DWE       	            :  out STD_LOGIC;  
READY     	            :  out STD_LOGIC;  
curr_state_debug	      :  out STD_LOGIC_VECTOR(3 downto 0);
counter_debug	         :  out STD_LOGIC_VECTOR(2 downto 0);
rst_int_debug	         :  out STD_LOGIC
);
end component;

component gtx_minipond_k7_ctle_agc_comp
generic(
  AGC_TIMER: integer range 0 to 4095 := 150
);
port (
	RST                  :  in  STD_LOGIC;          --RST low starts state machine
	DONE                 :  out  STD_LOGIC;        --DONE asserted when complete, deasserted with RST high
	DRDY                 :  in  STD_LOGIC;         --Connect to Channel DRP 
	DO                   :  in  STD_LOGIC_VECTOR(15 downto 0);    --Connect to Channel DRP 
	DCLK                 :  in  STD_LOGIC;         --Connect to same clk as Channel DRP DCLK
	DADDR                :  out  STD_LOGIC_VECTOR(8 downto 0); --Connect to Channel DRP
	DI                   :  out  STD_LOGIC_VECTOR(15 downto 0);   --Connect to Channel DRP
	DEN                  :  out  STD_LOGIC;         --Connect to Channel DRP
	DWE                  :  out  STD_LOGIC;         --Connect to Channel DRP
	RXMONITOR            :  in  STD_LOGIC_VECTOR(6 downto 0);			--Connect to RXMONITOR port
	RXMONITORSEL         :  out  STD_LOGIC_VECTOR(1 downto 0);	--Connect to RXMONITORSEL port
	curr_state           :  out  STD_LOGIC_VECTOR(3 downto 0);
	agc_railing          :  out  STD_LOGIC
);
end component;

component gtx_minipond_k7_agc_loop_fsm
generic(
  usr_clk : integer range 0 to 4095 :=150
);
port (
DCLK,reset,DRDY     : in std_logic;
D0                  : in STD_LOGIC_VECTOR(15 downto 0);
DI                  : out STD_LOGIC_VECTOR(15 downto 0);
holds               : out STD_LOGIC_VECTOR(3 downto 0);
DWE,DEN             : out std_logic;
DADDR               : out STD_LOGIC_VECTOR(8 downto 0);
kill                : out std_logic;
state               :  out STD_LOGIC_VECTOR(3 downto 0);
count_lock_out      :  out STD_LOGIC_VECTOR(31 downto 0);
lock0,lock1,lock2,lock3 : out std_logic
);
end component;

signal rst              : std_logic;
signal start_done       : std_logic;
signal done_pre         : std_logic;
signal lock_done        : std_logic;
signal ctle3_done       : std_logic;
signal en_b             : std_logic;

--DRP-related
signal daddr_starter    : std_logic_vector(8 downto 0);
signal den_starter      : std_logic;
signal dwe_starter      : std_logic;

signal daddr_lock       : std_logic_vector(8 downto 0);
signal den_lock         : std_logic;
signal dwe_lock         : std_logic;
signal di_lock          : std_logic_vector(15 downto 0);

signal daddr_ctle       : std_logic_vector(8 downto 0);
signal den_ctle         : std_logic;
signal dwe_ctle         : std_logic;
signal di_ctle          : std_logic_vector(15 downto 0);

signal holds            : std_logic_vector(3 downto 0);

signal rst_lock         : std_logic;
signal rst_ctle         : std_logic;
signal rst_ctle_b       : std_logic;
signal rst_ctle_pre     : std_logic;

signal lock_done_r      : std_logic;
signal lock_done_r2     : std_logic;

--Debug signals
signal lock_state       : std_logic_vector(3 downto 0);
signal lock_count       : std_logic_vector(31 downto 0);
signal lock0            : std_logic;
signal lock1            : std_logic;
signal lock2            : std_logic;
signal lock3            : std_logic;
signal starter_state    : std_logic_vector(3 downto 0);
signal starter_count    : std_logic_vector(2 downto 0);
signal starter_rst_int  : std_logic;
signal ctle_state       : std_logic_vector(3 downto 0);
signal lock_done_rise   : std_logic;
signal done_reg         : std_logic;

begin
------------------------------------------------------------/
rst  <= ((GTRXRESET or RXPMARESET or RXDFELPMRESET) and EN);    
en_b <= not(EN);
--assign rst_lock = ~start_done | en_b;
--assign rst_ctle = ~lock_done | ~CTLE3_COMP_EN | en_b;
rst_lock <= not(start_done);
rst_ctle_pre <= (not(lock_done) or not(CTLE3_COMP_EN));
rst_ctle <= not(rst_ctle_b);
done_pre <= ctle3_done when CTLE3_COMP_EN='1' else lock_done;
DONE <= done_reg;
done_reg <= (done_pre and start_done); --So that DONE goes low immediately after any of RESET's is asserted

--Start CTLE only after lock was just done. Don't want to start if user just asserted CTLE3_COMP_EN while lock_done already high.
rst_ctle_rise_sr_ff : FDCE 
generic map ( INIT => '0'
)
port map (
	 Q    => rst_ctle_b,
	 CLR  => rst_ctle_pre,
	 D    => '1',
	 CE   => lock_done_rise,
	 C    => DCLK
 );

process (DCLK)
begin
  if rising_edge(DCLK) then   
	lock_done_r <= lock_done;
	lock_done_r2 <= lock_done_r;
  end if; 
end process;

lock_done_rise <= (not(lock_done_r2) and lock_done_r);

DEBUG <=	lock_state(3 downto 0) & lock_count(31 downto 0) & lock0 & lock1 & lock2 & lock3 & starter_state(3 downto 0) & starter_count(2 downto 0) & starter_rst_int & ctle_state(3 downto 0) & rst_lock & rst_ctle;
AGCHOLD <= done_reg;
KLHOLD  <= done_reg;
KHHOLD  <= done_reg;

--When a block is not active, it will hold DADDR,DI,DEN,DWE low
DADDR <= (others => '0') when en_b='1' else (daddr_starter or daddr_lock or daddr_ctle);
DI    <= (others => '0') when en_b='1' else (di_lock or di_ctle);
DEN   <= '0' when en_b='1' else (den_starter or den_lock or den_ctle);
DWE   <= '0' when en_b='1' else (dwe_starter or dwe_lock or dwe_ctle);

----------------------------------------
----	Sequence of operation:
----	adapt_starter -> triggered by any of above resets to deassert then waits for DFE LPM reset to complete
----	agc_loop_fsm -> triggered by adapt_starter completion then waits for all loops to lock
----	ctle_agc_comp -> triggered by agc_loop_fsmm done and adjusts CTLE3 until AGC not railing or CTLE3 at max/min.
----------------------------------------
i_starter : gtx_minipond_k7_adapt_starter 
generic map (
	WAIT_CYC => 10
) 
port map (
	RST                  =>    rst,
	CLK                  =>    DCLK,
	DO                   =>    DO,
	DRDY                 =>    DRDY,
	DADDR                =>    daddr_starter,
	DEN                  =>    den_starter,
	DWE                  =>    dwe_starter,
	READY                =>    start_done,
	curr_state_debug     =>    starter_state(3 downto 0),
	counter_debug        =>    starter_count(2 downto 0),
	rst_int_debug        =>    starter_rst_int
);

i_lock : gtx_minipond_k7_agc_loop_fsm 
generic map (
  usr_clk => AGC_TIMER
) 
port map (
	DCLK           =>    DCLK,
	reset          =>    rst_lock,
	DRDY           =>    DRDY,
	D0             =>    DO,
	DI             =>    di_lock,
	DWE            =>    dwe_lock,
	DEN            =>    den_lock,
	DADDR          =>    daddr_lock,
	holds          =>    holds, --RXAGCHOLD,NC,KLHOLD,KHHOLD
	kill           =>    lock_done,
	state          =>    lock_state(3 downto 0),
	count_lock_out =>    lock_count(31 downto 0),
	lock0          =>    lock0,
	lock1          =>    lock1,
	lock2          =>    lock2,
	lock3          =>    lock3
);

i_ctle : gtx_minipond_k7_ctle_agc_comp 
generic map(
	AGC_TIMER  => AGC_TIMER
) 
port map(
	RST               =>    rst_ctle,          --RST low starts state machine
	DONE              =>    ctle3_done,        --DONE asserted when complete, deasserted with RST high
	DRDY              =>    DRDY,         --Connect to Channel DRP 
	DO                =>    DO,    --Connect to Channel DRP 
	DCLK              =>    DCLK,         --Connect to same clk as Channel DRP DCLK
	DADDR             =>    daddr_ctle, --Connect to Channel DRP
	DI                =>    di_ctle,   --Connect to Channel DRP
	DEN               =>    den_ctle,         --Connect to Channel DRP
	DWE               =>    dwe_ctle,         --Connect to Channel DRP
	RXMONITOR         =>    RXMONITOR,			--Connect to RXMONITOR port
	RXMONITORSEL      =>    RXMONITORSEL,	--Connect to RXMONITORSEL port
	curr_state        =>    ctle_state(3 downto 0),
   agc_railing       =>    OPEN
);

end Behavioral;

