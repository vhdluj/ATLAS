`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gT2RtN5Cdv0eO7GkVzDgI2oC6S3hOxxNOvy/bgAv6Blw4FwvwPuFz4XdWlFHnKSAZ8MBXntvn1FQ
uxyCTpzkvA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eSeqpNOKDnP0b2xJwBABi+bUSUh6MzRAUGA94SUoAU6e48ipc0OgExb6FrXTmLhHApUkIysdIU69
8ODj00qRqdzjHO2QHeHKPe04HJ63/d7IvkMi9zIbN9KUytG38w64L3zaA+h4AMzC6ymQmrLe+xvg
yEwxxtvrrPjOSgcdwvM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WvlyENOsRQDg1V15Tlo1CDal9vk+wffZWNilx6r39AOmqgo0hyHi7+BrnjTJrMKXpvihP+EqTlPV
2gE8ULcrBBTA3sxP+bD8qaUz3isisnhnmZcKn2FNdw7FLDfVy/U88MFd1D3aSapJMqEp0Il8XjFq
ckm3JmjXIzhVto7d7rav3uSO+NWIMsGTXUr5VJmK5+uYn2EfOSXgTuDJWYE+jkn/RFwtXOqDle9Y
Q+l8z1txvpxGTBtLp5TD0I9GuKz6g5Rjf41f/gu0p0dXyzp+ARy8dtg9jkzIXSM0fgnX0TD7QKf7
GQ4x3sw0I8YngmRiiCuTc6LcTPugOTL5dC1L0A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CF+y9dydOGqu/watDnYDkgWb5n+Jrd2W+wUSKKgA+ep5iDtN5Tbo0K2XB1G/oRXotnXxxJcwSX/m
YEEXf+Wo19zveyVSQf3i3i/qjc0M9n03iGKqlJXhUg2Ul4tdcX12As4QYueGL2zXPetgwQpywjBg
RnHn398LS33UQnIU0eY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KTgY7ONx8i7i6OKDNgMMAvSNZvdjiKfL83ZFXCjyhMVfq/ucwA+hJqw5jeyAn9xsRI47Erp4rIUV
R4dStYsRcPJGszcQSA1y4tFCanVkfR2ShqdDbBoJA3Gw5oFQeYCgaUqbsnCjNZxuCO1y1FwBMPxL
qmYw4PDAYXUp1fnWsCYaG5IPpdUnohNj0EaJuCbEZmJHudWN0GvOH7O19mBq1dXcuqdurZ5uvQW0
3xXvZb0m0YwUdbCeraRItJ04pXTKYtYeIg+/BRz0Kar/GK2OK2K95/oY922UHcumtEuYwlpd7ZAJ
JH6ShJtnv6otjv+M5Nu0Siuc0ZnkgSZArRCKgw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5664)
`protect data_block
JqF5oO211tf7tqkr9h7dSAQ2F98SorVUdjt17A6tfDUEW2y0J8tnt3npY1/1FzMVIX2Kft6aryWw
k9FZCXMoFPevvu50dqssYIzEkM5hRJhUUXoXU5CY+9GlgPjpE9UIsmAQKzsFEZPHLSyXQOfoKBVe
RWLFNetBVgab1AhPUMET8yF+rGC0W1oMs7P4ILVULhcm+zBynYKtcfJ8RDVyi03ehpDj6RoW0l7T
T9STa6ir/Qz6jCtRq9GQ45zUb308BrFvGUDmmoCiFFcsM6eBsdO1Du82hPEcxMs6L44BxJ/7gZud
kHiJoqLIu73iDtqqHLV/CqZZa0Ld9Fr+lS0yBdJYC9NyiVC62tA65eqZ74wPN46bIPJsnmzTwJsR
3DzircomN77iWNe0dVFOFBoTKpgWa4/vFyERgsLiiNRQQB+hxWr8qgLCNuXun+TDgT7uzrwzTjn0
uOwq6vJ4XaLLPN2Q8aX4TOJEwH/7w2E393sfaIN20SJsOw9Mn2cw8fii9d6wK5TZoG9Zt/sncU9n
/AuuM7Y5W1QzyMPu+tbaDIf7AyBMieou+8wSV03Ibn5XFfrcMkDWYnGx3aITKnagNSdMF7MpKhlr
GsMH9kqrYhun1JwuVyepbIWFNVBGSq5MSo26T/kru8I/zvD0zlDOZdXCobHDO/Sm1xb9fGBbF4CG
LdJIBLi5H0MFm4VZHOYHgFIHBhAu/Lu0QF7n61NioWnC0/jYrSX+pLgvaPVsznhYWsUI2QGKYfFf
xTHW8pnCUlIHZQCLG1V0RzR2lEWRQyBrG+cYZnAMsticR3ytZkz/zGHJUL/wccYOv85ZOCght6zP
CJtRpz7UN9N0n8EjyFOE7PDXUoFTnQh1P3sxiwhVLKWDJpLEzFn9eEtmac2XreWluHi3ISww6HOM
Ztcq0wZkcJjGraNKMAPd0Wnf+sW5OjPyEvUQoFgEZMdox2XBDQgBVOR65S3z/KKg1vRYi5YIeCEU
TVe4zxVvZIat1G/m8E8iIxnz8CwKGggSen0jjbZhIWYG0I+Eys47Gp+ruLykcR8OR5w7Cm8cTFi9
dnuyskvOk24K2eisg+MevkuMjBk/fLOFP4VfCZuRYG3k/GvPB2XLxYJz37z1YbBeYjuLLee+TQds
m1hJnjAQs4BO378+Jf3uRMEl6XF3zSfsEmQ5bERGJVO1QhB1BZ6GnWZrUSbFdJiECGzbBvYuVR5e
jloikM6QRHaUsqK5sl5Hz3yShfPqR2d2ZC8BGbeF3ICsU1JPXV8t+MzpHloOdA1p7lfpbfi0MFL2
yV659b5cvOp9lfrJs0/jp9QdwSGarXSpArrYWvB6zTTUYkBXlLx5hgUPe666nHMX87XCKOydtLzW
fVeRlfKdBUnElH/Mmb955Od5KPM4/t8vihaHhE4l+o0EnbDVF472bF7HvPFoeaqXDDMBZiIKLa0m
l8oJlGj/Ej1IqO/8p9sn9N7a1r+8Z9wy7mr0tYZuO73E9LdACElJM7pE22hzdfG7YxM2KMxLCjzb
tDsafA47zeFBE8JzZXdimpWoX09Q3z/ty0F633JSY2/mZK3inL6bpzL0xsXj1d+/sYIqDUp6Bva6
+SYOlMSgpWLI/yUkIZecprOc/zNcb/QASS8Q9S9yhCtGE3mRQoTwo57lQfhTsu/ioUrp0ZISLdgP
rjQ8r0c1BSF7CP8d/8JuSfiTuSCpn1rnTBA3oKpNJU4FvJ0XWQRbWNRNtOSqzGLxFcykB21rKguG
1jA3qv3SuT9QoStCqH0G2zahUQypSX3iR+yqiYCsWPoRxYhMCDgM5oopL6kmb3V7SbDLtQVYleoq
ndBZRLzmoTuvqkV9v0agL2E3vVGdviFjPgWnZHN6TdU/V6UGUQsryb94VolRRWjM859mXNcGErzD
LXTO4t5n9IGj5qT6fjwO9MEsuwnrNWmgHFRgGtqC5wNB4Noq15vFwkErgE0/oS0vfCmLiXpuR41x
o2Wf6GS+rED5iMI83mVJwW5taT2gJNYslqntf5ha8R6fB884F8N1c3nvtk4aFBz6RK3AXaHh75Ty
2UbPhRDLyvs/NMnjKBKXjArpWXqf49ADm8qPaUZLfPP68DzxLkAR/EPC9EHLvvQb83eHFXv86SlZ
u+A/Srou4a9ezjhlsew0nZK5q0PxT0qrhDP/1nLsGC9DY/vMm/kOMgtTsPrir9yubVsAZOG5d8Rv
OM8xCrgN0A42Xh0uNUxCgjyC5lVn2FJME6KJgaSBfdCYHKsh1DlA0HO9Y1QqJn1hY0AWglNuB/ii
oksnwgsH4aTpFl4qpVMPX+pEwCdZl78ME31R0VCf4bop0ZjI+w8qgUBwPPhnmsy91A5zHuNmqNIh
g6wj2TPMQg7Gk+MXHtgRor6Nml4Kkk9/HzR975ke+yLckljX6Q4hRf2RZym98lBQR1gMdiSskZXz
zCmQI8e7MXVyljk2uPcL16HxgEblAXl94ZotQ2R8QT6x9pQYjDfWVN4jEPl4mMq3Zt0s1+HsEFhm
mCVjlbxqEvmQvw08mK3zIbGYnyU76cFEu1UGAyK7jGlcMlxZnD0fsOTQdPMTZvipSuyZi1hSA/6B
lL+2BtrxR0AKVRsb2aBEwKwFBlONHQSD9DhJnD3TEW8R/tisEM8UHba4Gl8YkL0syqVH0Yy2T76I
veZGKiNQp0AQK4MrltJoxQPuzPnywmmhkLyljIFHwEIAsmcnQmhEpBUKh+9mErzyKwoCb1DMlpuz
RSFVLjuBKxBrqTRLgqUw0HxaSrqoyKH5VmbtiCEhpNmlh+sB1+74SQLuVfdrZKD0B11ijM/ZJcco
a7GwvdoWif3iYb2e92Ey0WRIxi5cuovE3yhOcKA/h+QWBiAnP3ttLamgaTl6kf8gNp+IpcDCPJTU
/d6fOc51a+LdawQzNf7PC/KbhHVaiV1seLZ3103kslWvvLancoaoN9bHwsp7/4asas7v1VjsBsQ8
qzLUqU61yA8idie2JZvHpnWfBpZZOJi/SipPY8zpPtMF9hfaAL/d4NzTAIwHSnpa4iG1+1v5MCsc
yT6azb6pSLhMkF3PJsKG88B7s4PCZhliZBDpKZfj43nENj16JCZuILAPvctL8LD6G9+CtSTaxO8d
3FWrHNchqkcUm5vIJ7zAlRao9sXdcpp/CGMJFFydnmeZEJPy33FPCrTbwpSqlqwuWgZmDr/6oC0+
6j9V+9dxhtdMlS0Q/tkbkZG8rIjdt/XB/gOSyo+bGMVCS+P2hOEiNrUH0I17CI8QuZyUJMQtN59V
WPAkzMkHF5Wzz/M7oO8TfUclc46ZmIQW8GpriIZ/jPASScIrreeeirJw8OIhncf9Z9K2CA/aES54
yl19XHQoxOZePYOs+LS0tCK5BwglUaf33jrSM3CODM2UebfMGbE/oHKdePY2kRGp1/EPCsIdgMRM
WXxtmRP4zW03YqDvO23MxC4E2E0Jrk/hUPcu9gajG3l9A8MZVg8TXU/qykCMJD6ESWsgTZYPm0k5
SYD9NJcd9F/Ybn4Dkj/0sjkX6faZdoAFT2ZEmMhxXsvgsbvWcASBkKEzuTAVNDpSfH3zSs1qyR8V
Ca3wdMVbZHNa3+S2k1nqXHvvnsk6obQhc2S8tK3p9IVqGpHrH8z9jy8L9TAu5kIYG+GogMCQ2eSJ
XLTHEbJfvBQX3Wv8AAAR22z1B9z3VOBZul1a2KCQTKkUDKCcCtstRylbsSOz7Qni7HhNyy/HQDuT
oz9e10cK5TYXrDa6CpFYt5p9vNTUgYXgUvcUgTgwwLQ0u3S+nMl0l6dzEBOA0h7a9G60jMFXb2R3
J0KzqIBdUTyYB47aWv9rDemVzs6YED6y50WdkGNy1f6Kuc47Eb9B277ZbIHHBtKBePcivutoumMe
ZmIIc7DoijuagNR/c0eQXNBdSxrTVgsAzvXhupdAJIWr4+AdaZAcLzIMqiRbfRr00DXti6VvCu5A
CNWYQeIG/QPxtktzOO/+Fp74Uj9iauNvMFdbvwPGTDSCA3+Scv9d0k5cIxzB9KisePQyR+t56G/I
mMtgFd0EWrTfWOS+IcKPZp/8Bnk6h2ijB8tgM43rf3K5uIhWt7qhx+/BGo2lxH/r45LTe3Zbr14h
mtvNStrKPFQ0aFvw5ajpwbzDcu70dJRTvxSG7Vy63zf/rve5/vg0Rt97gb686Vw7b+bEMTeWaqLu
x7VAtfcLeFRSDL+W4P9aD+E7yJCNEfvNdQ1jLxISNXGziTZogSgok232rNdAV/g5s+fSisLsDh7n
TYD9znH0fRq2L7q2jbCLdRMlE1TapZHd9upeSuMI397sEcs0Qw360gUn6hZdufZJP7OFMOmIgUV3
LXaTB+u6zY2HkwO6CVyzqqu200sNXexY2aWAHKfgzHv4v11/pF1L3PT72qB/cv4O1VNqaHR34k8Q
4rnUBEylM7t+o337w27Wpr982qQkx9AdV1zrorm2EvHnX/oaYVXhAmPyLFNqYjTSg+BtjFSBQsvA
VNBRV3ofeB6msSO9BND6m7HJJPHhxogTg0Hd0VVeeyJYU6SLKSIHgiG+3fgv3zUYxcm9NJgwwMuM
ja7F66xhQkvtvqBp2rFSdfC7XIeattNUOkf02psAcqhPaKjshZJfKdLXIBHaU0Fo8ucTcCL6IFmF
NkVriaFxlyunV331Ae4IGnOZxwLU642NwU12TnX6jI9lvp+XP509LlplnLFpu/Udhpbu7TkbI09i
4HZpyjU50oMPGWcXv8stV83rw3rjfp3sN1psxHosM8Q51OzkwDZwYrtxPJIhs6FoiPblTHRu9WWH
44cYhF5mH/IJbetrd1wO94tuGD54m0oNqOe2Lxws/UP4rPE+QptJd9EIYT/KZSJj6JL3NaR9Ys9g
cJ0xb0z9z5V+5HbmGbmSDJxbAFM9h6OEI01IdHnfVNfQzGDdsMJ2LDgDaYn0Xld38RlLzxHXFfDp
qUGUiVLUy7paNZQmZmDqQVCZzNq7U1Pb3nUUmrasHkC0JIt1FdhsDAVactxSPJlm0pa26cjazZ68
vl+L9ViMkeJelyWU3lrTrhZMvLMzc0Fy0gHYQv8T/nCdMdefool6SpMVgayTUwcFVZKkbTgTyj9V
wQMlLztbvnOOmtYJnPiHjaIOe1ixt/k/0hHJ+ssZ9XqmlVa3XqBo7cB1AQTzMyrnQJjK6Ro6+tLy
65+EFLx3sqirMxVP0FAPEnXiPimWhuF7OHCXJZOMhM0bYoP5B/0u90LP1bpNTQ9kdZg3UEXQWg3u
epTEnYcfcSbgaaNYPERv/fJkB6tCwFeUlU9MwHAnQFqhZbwiEiLw88n/sK3SRQfZVPHtVsOirC8+
TwTCWmHQLxCopJKjMGdapEZbrjOzb7aXtpVAaAQE5p+6GTSOnzpXqCgXxV6B8VV0efsZrCGXhNRX
cpLOedu8T2T2S6QbWcoGTyr5cUlTlIeOCGTx7/xDbJ2EI76/kurZyg7u/2P7u1BJKb61JDvbMC5c
GL+9AnVwqj+lZb/50N/3I+NkFAFJwHc/9xDij1UnbEYkUw8e2LifDp6lHtsf4wD00ovbbNSN/2pr
D2c2r0Xng44hFHrmkNHvgUYecpoQSgruJeuxjrGs7df6W49DhiR3RNiNIbrGzkdY8bs8NeEJDsSW
fV2XSdd9xX8YfA3G7xf0gVty95NEbdsXcbX4jo88UCvbn22o1S/oxH3TsdfkTd4flGQZSNRoL4Yi
C7qClyT6jmV1CGhhxL2CTAJU+im1McRyeUt1CQaLjNDzfO/MMA7kEePJwbCKDk24KK/IWF/8AGd+
YincmQ1KqwjJwmeV7n4loX6kLbRrzutt0Wgquz0zuBzQvFIB+N773epn7S6KOYL+gS9Ee7l+fRzN
ZAkYs04V+Rq7aXOTYJmeOOH4VMv4zn9WnL0gvJftlRyA7HTN025py8uUJa8x/MuTCNA9YplcKJhJ
+Q5BR4IlcuItS5Xr5ZcQlF25SoqRZ3AIoQGoffGzu9DjxilqwmYpXJAgCc4qaPHknDwaT2HJKJIZ
tGms8yPxEHkqN2MeKNkb2FT6Zdc4aMVuj5lXfr1p8VjOJh+UKGOvxU8K3TuxRcUHIXD9BfFFHLBO
yQQyXCrgH4P05ZCmSql98/pfaecf7Saz56nlvIkit5aWqNjg+9TRxkhbgNotpoLL3AKoqiXyfkz3
mn+i+/6zUON1N4+fU7eVKnz1qokA4SB3/kuGW7elTDB3q5fum+KqH39vlJ14z6H9GBqgv5ZFkAjV
2311ovJdRz/qOvd8gFkbxfmNNGIwfBXFdYoF0GqHlt4bZHkXYxpiKIWF1v++UElvHSB9ORIsgUtw
h9AET+ShokRybwIBhpiBq68zzTdmxnQcGOvjDv6ojR6+1qG8n6/qvuPWO/4XmaVNfuoPaTPBo3lI
WREiOUO2yPdQnHSsj9Rdp83TQZSIUbHBc8NL40tMunUSSasqt6ACRPbRxcQSbHfGF+y6wnoCy9Ie
T+wzwRONmGEaXooyvMlfFiu4KMx0wa/PkizAKI6bIzUDvCA3N2iHIscPKQJp1iu6taiogEYeIc+N
Mk124iYadY49LayxJR3fh1neMBddGYucBEvoGtklShu/7rKaLABShi0IH8LUckhQqvHz6R8uO9D8
gwAitbv3Ji99m7wncLas9kMR0SrauAu7mLWauizHyq/CsUpH9QD5xtyMZ1NH71Xf+dfNsRSnULtZ
Um8HxBGSnwERqScwMn6i7XZs0CFIvdLqsUD3SOe5/xUQfA9BBi2W1q7invuBG6OwYxquNTruVNFK
leppQ0pvsm08KVQ2R8949U4Ft7yL5DMaJ8Pxg5lfrzPbmovsh6IbmGwXz7fRXzJDP+EcQZhaWq8J
pTDQhpXGrzI7ZrLkUGE1TTRs+trYWCpDdpn9ndWbAHqFFkyV6DBfQjalWG/EZApDA5/eyz2mNLwl
KYIXeceyNmjMC+4c1fXHODNxq8yAqR3Wqx78A1hykHUdfLqkQs69WaB1NKK13LSXRHKug1n0bgH3
0xLColYXNJTUv49ftnN5cZqe5kCKhqDbhAkzt3eeRmKXFJ8eGHKzTW1Stul1OCLZE3hZjox6cbm1
PwMusmfL04sgHCOiDrXGhkjrIZD2Fuedww3LOKa76ywfUcPtwxC8ZpOaM0waGjF67RlMuK8e0coF
8EuOPorRx1xGFOkFGP8VF8tn2jw9rWDf8jk+U0JcvoikIR2M6bVN7Kb2RIp345CB7xucpu/BxiIi
vQDFXhVOjGGSFAdJHVmDZstqQRlyb6BTJkTUTyX3u9HURb2p/GdyjUFrNGtqYhneh2eyd8kiYOJE
znQ535rE6Q1VhMTwN9Y7b/26sFYV70BBerdnvwlBbDZgSDh9fV2Pju1oi9WsLxilaYy5OWQkBBa4
xhRz1/DWbzl2DcnH3AwQCSYhPOn4HdQTt26IAyTMBJE8kXOJdutLp8xxutcCmNm1eOzYLPAYf05n
VPmAxSJa4V9YFLEjBtJogmFEXJ/2Azd5no86zxjQhk2ngrtVye9UDJ5YmDFCivm7PYJ9qRC/Km96
oWg9nqvfudqr3mF7uFIJeX6Alsoj
`protect end_protected
