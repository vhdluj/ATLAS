`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BYcBUY3bxptKfznTjVHp66RcUUDZKeCY1jthH3XfH+mgv1fD6VH+M66usblDc36tzO1ZpWRaO+gR
h1IdDcns7w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
paVNjPJJYOcFD0smHohPi+ia8khraNV0aF0BYYlHeh/IYI+hP8N90XcC52uirU2VRDXggOkHmx8s
ju8kVgqb6Ty7Wg22SiTODknToLaFY+K1ZT5D0iKRE8S01BcZh1f9OfbkiO+ttzozes53DtNvP9t1
5eHJrN3jzaqqh+rLrpg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wWUfNDveAX6heYMe84P6eMplyJHc8xSb+AHd1FqwTmJ+oeme8RI2sQgnHNrk8p3e9/zk6S36ZZS3
lLYRKXsE7Rl2KzAsfrB0qkhMPLK1X88+9eOUpk+Wnm/NzChVNGLxwbItxvuFOAXs5kYOZ9H07YzD
7b+0SLnGB33wLxCqvx7xBLQtZr5UMrWZ41jftMa9PK6aPdRBPHisg8FkXs/pS1mjCtNnEImijpQq
fHl0rDKh2ts+ramItlMeJfqLvFgECbhR+6/piYDtuTkBltvH24Ty93H/7RGY4I7wzuwNIiuGmNmn
1aQwMsSEfagsIi3+zeJ0TiKtaDMdF5oTe17nJA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3KBcRf2HoPt1esFrjs2yIzaXiVzykH2PB8eq7maKeRmccm9MWAlx+COUcZRCVdxvfZndjDCGzWNw
WCJR+So/q27udrTm6lI3oy89cPKeuxHlp38oOh/Qfo2z1mYoZ5KrcxBq+U6G/m6Z6S4NqbY+84x0
m1B1+BI6QSxXjQrANno=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rxPBB425FwLnZd6+C6ZTlCfr/lqbVbqMNyrRbeZU60d73R7G8p//ek39b61rOG6eRYq5C0+sdb51
ef30IRakI9IPoS8zyHgdjSOc11zwHFD4s40B2+rnz6w2BJeXkbVradTuXM2yCyGjKwmMnb9qS6Ay
TF0RHNt6jm7J+6N7qBzLvA+zMNvS8+CR+H9oCGhSy2CByxRewYbM5jpzwCnlpF/qslUIgzGCdC6i
esFVq0ecsJtMSpWlLHuElMf4vxcg3pwtn4hqHcPUXqCd7IYOXvhU467CLhTqcJDgthqYPcARNO6r
UZl4p288j3qnkDJl2GFfRGCaYkCJ7J2g62HIDQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10768)
`protect data_block
LoExJQGww6499xwouvhcILUr5N8t9xE/UggZlYDoWkyfgBmP2TikpEIjO3QDK6iFS08SwMlVPpXp
fqFCRpQXJGKTNqKvH7HSqwmFc6dm0UmbEwcSlxBla22uctZmVUG91TRHlQ+uDTetnI+iPqzv9azF
Kdf43CcuX2ExSzR7ujNoojIvQvApQ/GhIxXodxwzqr+5c3sZr80uuqDJ9VS4lXNo1VZ/cesQpGMf
GOiKodHchn3UI7oKrqY8YE08x7oJW60aCj8oiimx+0UZsp0rI5L8Vswke8oRdA+gXtybVuo82qa+
TIDhuCW1Tu5gfZBi2de7rY4raC4zzMJw7VtSrX1QXTBMFRAjOVTlVGPHUIsfPVdmx57FRV41kQyN
HNgLJMEqH98jm4M2BSCGBsOECW+bwwmBMaO7VTxKN4eHgvIbbbE9dQMlXezXEVUdupfMr2eme5tk
wChiiiUfyc6C9f8RhXcot2gav8iP0R0VlQ0yXhbycKV7dihKwtJCIVqoKYn0Mh25eSN8e4jWGN2D
qjOT95Zs7vUIQtgR8iCZkzzRWxfIU6fEWEKScVC7Qhu5oYg/EVawyznb4JAlRjb9UwhxT3wmuEAn
VxjvAcmfcSsseWvOW/cXSDG+vTB+Uk3k0CHqZLoYlmQ8KEqicmwgXV3zMwC/hVkcU1J5P8UGXExO
GODAXUzGV2nF8w113xB+GfCGRoZi6BY8PjkW09F926tD0mK0xiL6Eltb/cEr4XcmlvJBXTukcLVA
248UMdNNo//wnvj2aI52hip9ipmgFyOoIXaJqgSy+ahEa70en0R531W11RrLU6Vgo3PmLvPX3JxB
HYdPUCzLHJCd0E1QB9drWx9nXLA1gM+IBTAWc21KwVlnP3jSYkadk0m0tUFLw2o70Iqc6k7WwXa1
6bZ+KwWfExpEePTBkmSDEjdlYWo4HCh5sBUKRNZ466ipMVF3smSH5Su6cDqPQaKNVtH/rl/kB3Bc
tPpaG8kNTi3+eNFEdNeFtDOFDH5A6GziUtLYsjAq/fTXqnPLyDyZKGU0WeCS8vbfNdkvLFzSTToz
Gk+LlBCs/maQevTLKfIA8U04Prw+vz5nn926UmgY9RL+5hkYg1pW0+OCApmKDLq2Zx6NRswKCwKi
Uz/hSeGYRhd5ptEziiVqtWAtokJjQj6uFqOxBtxm7R8xOakiAmx8+2sXTgN12m6Ttb+1a2Y2/cmS
R09e9c8XmdKWrpm853JuWq7OHG7SFc5VH1//w9AYBZjfxiKOWQdIil4DOViJcoYFtlkNNs9vuH++
/deVabHE7bLTiG/6JWlqeDfGOWS+2ojmzYbJEi5fnX0v40mOP4zpPf7BFTlu+RwbxztHZ4QVHhT/
B31EC+gml7/ZdGqehGmW4MbLFmDmxiY1LuA7OQgu0RfXQ/VfiJuL1GzDF/05Bnxelc821S8ctf4O
yxjiZQH4CfYrdGLXNyb2ZPeVxwdwAY0X//hAZEDHxkLpoiIRlwtH11tX6o9q7HNSCewnO5wOa01d
5fRQJqy6PHcHboWggeAAC6udyBLJUzSgoOJwg/GGQ5D3ge7wGrQ6HAtMtOszaUeci+Zo4pkoZGEa
72VI8ESSYQBO7ZHl+KTd4D3VS+Qye84QxIi0KI3H3mj0oe0c6QnqHq1YXjKvZRcSYJTVAUg8aAZY
QSFVT930dQzPQg/YPBZGdp1DX9ya1QvI6XjKPGqjWtwPeK5CjHRtEIU/wrwA/4gkPDVtuJY7aBdM
kqcC1Fhtxy8mqH6lL+FZfqVmamWKSEzO5s2D5ifl/r/hqmpw1orugqoGW2U3MvtKFRZQx9lUgz1v
ncEBkaLrWPkaX9IgMresIAIO8rCLiPtKuL0CYy1ckcQbkWR3YuCZZxY5hpJZSdpffJQ198E7dql7
Zv+WJXmyL89Mk3cjVXf9UuvDKzMb+Nd1iMTOXbcEgb4cyDQXKkV9lOBdKtu5kykn9PHlpFLkc/cL
ZfThRIJZsGgaJ5r5mJ/vioU0cLQrnW8T30mpYVT/DbErT6CbarBKmaK2vwwr9ec0AzZlR734gzvJ
eLFEWnSRR2TkW9Kf+twDJQk50XxJ5AQFzCX7w7TMboAKVeYIcbWfXThFtIa5gCTaiV0QqUxEY1CL
v01kaMfr+z+cfUu5dJwn0CHjEvK2p8wIJ8dQD9MISerEvR4vd4LgYxG2RfgAKBwjTenzi2xXi0mw
KMRjbQebYGqCG7XAryxKgYtoXWOgWwDzm3RywMx+mLsLfIk2WbT8jOoOqJwNJ22dPXk4lqZ8NhbG
QEuS+lVIMncKeFP5RyZJ/nFYZwuBYwT2XBEpXseCF1wTD+uTV1dvtVdwMaZGEm5qYWn3L9jaJbqm
P1n1pE2vUJQVlq04y4e83X4pnvLcwbn3wVMdGfCoYjmFDvcvBwctioRjkUHfDpXQGR3U31Syy+xa
z6GuAyyR/5TXsSGfDduwGRPm4lo46LLsIKQ7iYJldwdMcvOEeUNB5523SwOABgihGKAv82u5uPxt
IWfzVUosaedPKa/STZMpac6z/KWYPr2Da8kAMmD39zzw0ZRjS2VondLzW01UGz3CcQJkunengi6R
nxdac6ayS2MugdtR6S26YoPmLzWLoP9eByqJvH/K9Kma86+jLYYKAs24Bb3bZps+qmZG9z23LZDN
zYoxcli2isNDI4ImRFofrDyKcGJz07NgEBBZCbyjvTSvZ4fAp/P1SkS6lMENTOvnvujUFvLd6b2d
f6cdp8Y4xhGpZTCcgJ80/+bh1pVdh0NKhxDd0isJCmAKseYcnhNuvL3VqwGu4+F8DaQEetjQv32C
Badkro0XxLVwvVSwnZ/hfl6hrFX08hCYhzB4N48FwHwE3pUOqjeBJvrqm0fw/GY8GVMhjXSDLGdb
vC+Yqh1tW0iHtOr3xOAbf6yoGAOmVUhGEjJClXBetdvASxkzfrfIgmfNLRKq8eLxFDHWAhk0q6Xb
gtd+ElIPARoUuKmNLAxHKgO05Csc7qn8G7X4vBYnJybac8vtvbBA/88a2BfmK8LOY05W2eGqx/uQ
XqvXI1w2HoqO3lQhnpUyW0TWZfcriyZUGvlNnc5TRvLSTY/A1yKi6B/F14e3YCCi4AOgl7BmRoD0
YAfqYga0jPkkc5v+biIUpAxpTOAv5rJKanZbzHPbetwTybJtwgMinAyuCoaE6jVI9+R/RQLfkZzm
E4+5MntiBIzu2QqyRwrXjKWwPsA/4fBnlVWCOg7lbo9pFtiCR5QITqvPnT6Kv849OUUfGJuE/nfS
0+zMiJDVkk3HgfKC/KjVjyLLV249dvOe148wsROwJtv7HKcpv2+7Wlk10Lu8F8Rf6RFBQT9JIvth
8rOz5jap7gCuA0UZSclzB1pFAYcqkARjVUjc/yzLxG44XE5tq/g9zG9JOE9B85HEAtgyqjpOw2Kk
J8V7lfTEN9INa9NsSMrdmdJpAoeUgk6/8P+mpe+Rhfn7/GJRnh0JxBA2U3Zc7mpfxvVpGgSA7Prh
lfLOj0Y4lgDfx6F+5NQ2z6mS+LzEHSNfLxKXivdIVHDeQVCqonExIIoFuHKc8Ud999NGiTYYbmIs
2Wn97Izd79Noa3SerUoHMB0ewB0kGKhc7u8Xj9wO+UWz+p3ZhFUPjOQqu3P5NKNEpim/MCzs2MAg
6iVT4GeBfQHVI97UzoD9LC3g3e0yIHDWvz2FN60CgZHR2k/fHisAFfHSX7c/yV1yh+yKZxQ2WriL
CaqxvdgC6oW9hHUWD538C2icrssbMRGCXAv19lngkRlJdKbMLGGIGLaFjw1U4BYgpd1DBt4J0KRb
HfWOhBY6W91ndVjKLwCKh6elWgneCXu4/km+vdCRI6Uxy0Fnu8N1Vt/91nSybJUSAp7/QJAmjUkB
2GjsTAbHOhGdjlS8HDLpAJQAKk+Ph3iNqBBhPbrBKqPyuFG1K4lVdXJ/9E2CKH6oNqWFx8PBUml1
MSlnnA9QH4jbt6CQZxo4T3DM2qtlE5aUSOmRvfrHp7BKe35rWt8vdfdxDkqABiqoVJNGgwRnuMjH
+TH69b11dWaqMIAWW1idBR5vMvnLtva+tfeRYsYJi5lrzqJFoftySyhHpQNk3RLzxV6pGc6vwd6I
TvCxOL4gkxzTIq4mD9JCXcAdlk2mqVRVby1aVoFm4pP4arNZrFFW85ZnK6FS8B8SAM32SXQwrK3g
aLSgYIz18k2C3Jb8sY2aZvtcPlvtn4aTDaSELds97M4GmB9zf2BA75uxTSuf9XwhQjzYb/JnhF/s
aXXOvALA2OOr2Rwl63jzlnkOjfwPmihurKDcwKpSbkicZYa54mLO/Nh1rMd4u3aLewJ+eZOMEp4J
2NDQUKSvT6gpJrGWsfk6jl65QSPOadzlGDALUllFpUbGWmqludfbiJButBEqTR/MniRqhp4suEHZ
JQUMHgG++kCtnC/DzosdyHMiEgVj9N1puiN6OUbIwlZdtQzEhU96LrEf/aUfejR7ptd6wfIYXQrI
22nOtBGnYJCVpx5hnG79ADw2yUFFGJjzR6XwWUCAronMXQJ96ZbOx0sOTYBTpEDearTeVhKMdJzk
0Jaav9Gny1n2LzoYesJfqF2+2cizrRPn8pVvvJIUQiO4X5C/H3aESadJBr93OAkEo9wJDVy1oIch
CVtpQpAo3trDmkSGdkP85CXNcHjxdLfZ+trP3PRBzdH3GqQqRFOvftZi64dkG6hk2Cp2ZdfB5U6o
otyBVHjAsdyegLbkyGOFHHof7XpIWP+yShJSoMhho4GFW+lQFEktBUbKfAYyl8lUkdXpbU+ejhCy
2eQRZmY5tU4eXErccTrTJ+MdHBo9IPae+Zn9kWjniAo+U4v7Mq79/q7f4s0O6jlNIvsNskFaWB7W
3Ay33kxIrRnWQv/LXY5Q/GxHMmPBZi1xRV9EcY0ZaINs1+nsWIvMX7RuQMIA8ESutkVVO0PRk4lT
yQ+FYjNCbvaUpjcX2DoA9hvUb9UcPUv2IChZZEqHAIc5bcqjIccaYJk4tGXUlT8Wfq/KgxjIVMS1
csxvzOxpDmyccqUXT5FZ+8wmAooW3mdZLCkE/jKqdb9WMIcDOUqmTdKQvo4XHIZ0AE1JeQjMf6QX
rOUT54gHVqj2zRzfDXKKY1ejRSiSjDkeuR1XYNsDnnHO7dqP6S7OHhyqhPEjAn4suBkcoMRGwO0j
IoHc0Q6UShIdhKBhE3sqvEKjApbpiKL1MXW6qRCnz2PC/mCMjia90IG9zjpCPloQPZ0Y9mTLuW0E
hxMKHKi6hoSr9MXQIAI9L9wFKpq3gY9/DlwUbMK2Vya7ajUu8OjiawOs3Pfd8P+BfYCBIrsvYLer
a+mu0ccl5ffi9ING/nYljSs4wdvig1/jXpi/4IhXrwy5xD57nOTefpCEvK1ZIKHUUJLaOq6l12iL
qvyRHL84PnAutKhX1K1SxyJFCisQ5rnatMtDZiEGWkU4oXSKCqa8GUie/wii1y6KAZlqsxc3kI+R
Ky3MPLxQ62VclfgusGXTG+fptmOFT4El8XaMxzkM2Irba3eYGiwzw8rb+OdjcToRLq7SpafsVuIl
VKMNTPuRJLDSvIAiW2o+JepgWb1hb3DlnzDXkNbYAt4Np8ptJ3lJw/L9HFWuFcxiz8oXtuxYrhs3
vokU5hvquWu4nvK6AjG5RCPqONTkhAZZgelIfUHTTMwvhVk9ONqYWDOMoE/WZLKbWunNvvqH2Lg+
6nBABnpLZe5YVYgft4AhAyRs+N9h3U3PTan5BG/GWxlkJqnfK22Wn9I4XyZ2VsS5fEU59V+ZktF/
ZSYEGdygrpRczzmtB3N30p0uz1tpYhhb8W/9dop8Gir7WGI+yJjmfop/qzVxTShGnhR0pRoGEYFc
uGz5SnBt6WWisMLyOlkOgvlfRiRtBBFRYlZn+24yfoX9m0g08gY85KOJM0ZYcc6y+QIyBK66TtwJ
kRiwty0MMFsynCHBqtVOof4ilJV/CU3szLs/9YlvHv7ok31upGt3Kf75+GUKT8U/58yNQqlEvcZR
fZ6uSYCMD9mkirjMgzuaqn0tEUupY+n1QttpBw1VDbDGzYnH8dPV6w7H7zYGMJ5QMpo8BSw2WrEp
+ZZznvt3xduMPvKuBUaQn96+tDZYada0+WVH7Rx9dL4cDfeNwsYJO05mlWd73eWu2aV7vZrpxVvs
KC8sGc3dgK6fdzhr8BhnPjpLeq/C4Edf975SdLaRwFwMUFIjBfXF6SlJ3Zcu3qiOwy+ZTlAMWKAn
uf3pJMlvzPKoOfjZWIxiPcbseG+BZRyiIM/+zwszsYH/ucy49l7/RdnBIyQOTHDzGWDHkL2XgL6x
cZReq0LyORsflAcjpvREW8Q7FGl/hfkpaqyTscY56U4J/0dHa/PO6jwAIGHvoNCUIXUjgbT2zV2o
mzPcxcGSTkzx0ZAE7iit9H5IwQbQ/vAvUdIDTKqd8f0pzSxw7CZref01Vo57bhYeav+Y+ruMEkuC
MBXHqrB1I+U+C/HyWudvmK2FARpR67fGUQLmxPhDWzzJfLXPQvXh9SzueFIzWafEPm4bSS54AwOu
spIwyMjgmsmkwSONp1FVNpTA2EAcI1otXkVJA8YAeXRYuxbq+pQrrEiygpWc7Ndr8uoMu+jrqxgW
6q/Ty7RTuov87tDP8k+uoUkR8I5s7DE35eabH7U+2ElrIQ0qnd7FboO3MGpRvgl1gXQ/9b2ap+m1
ZZrwDGSfsv55RA8NcEu1eCB89DMiHTwL31EhWN72iAw+/RVY0aukwGPhOHYt+4HToAQTAe967nnY
7MPwa5sedQ52QMhxqahnaY1XlZMjW2sskEJsIVRkTIK7p/R2kPR7/42cP0Usi1bPa+VrBsHoBt7I
zAsL+ImU9a0qpjOLVSGrLNcrpbKxBD7bVUJQNIp2QGWkFiCgZw5GXa1stMf4Yk5/4pOocwtH1xWi
Ghi39pqCsc5mqPF/rG/RqZlewjvmuqr7QeUKFCfZs9Vwjh6ftjEBv3BIPS0BiLss9T89k/zujxEF
8qZ/k296M/h44e3zALZ0OdSS5zi2tn8/ZUORR4gN0Of9YJTChenJKyVPsDJM0BTe23M/7YjYOtb+
pWfOykKvidddAPF/emourkCZC56amSGrUOXdICr1mitfNnAFwI2yuw7ThVVVsqlvlt9Smbe60OLP
GOlp6SwCQ5HeRzP8Te/RCFJYWWqw+qdoRU1X/fKBVqp5u1gHb2F2DHUoLX7cIhnnCr5LqaXa26lv
uBwNy8G2zzRv9aRhj9N/3EbyhNlLjMZTjoT6Z+2H6UDKEFMWwVi1NspmU1sffAXKtx149fQwSyd6
+H2syE9drnUUZowI9dPe8Df6Wp+y57FeGNqx29pFbjYlOck8v2nrXPbeSfNIyhXvdN62FIynHb4A
0kozNJ6Hti+JO7/fYy1KkP3jscB3bWCMtqr9nHNj9bQxaUAqgFj2D3VnMY3PeNTZZpSm5y6IIuVY
2A2rfV9PJN+jAR7QG+iXVzrdPSzAUkZRvy3Cu/H3L4eDRIZ5gdWxV7Jp4rY9QGQst8YLVcz7LSiP
q212B8A3SunSaJ7A+hB3DIjp4NQp23tq6AIXYuNk8vAzKNqOU6Iv7poy657Do/Q9Q/lisjNK+jOu
on5WMXvgDNbd1RfvkRn/PreghGigQYmIyrar6Y0WGzipg6vMRlKt33QXO8XwpbqMP7Lh4lWBkvlQ
y6bu1MVrID9kM5iABBNO/0dj3qUDDr1dQRlSM4lqX9Gwudo3b6Bh0pF+XscjOV7bl7PugvHMNBqR
s9fKxzN/LbFp+tfAKH+jMA35fS2z49SQB7YASkcozD4v5x8IRPHNTnzVH+sAJKvpcvebqwxid3xx
XRe+dQNp3bIUoL3h6ulZ5Z663Z/TowNhiqDcWMC0fmaN9aBCal07bPMjBztAB26dk5H8FqgqAKhl
PNMNFbxqjBir8rOQ9wV0A2NSOl8PiKzU5V+GjR4SE+nukGgLuhTocZ2cZC/i5c9fOradrqDu5Lzq
GLg7I8pp6MsU/+WQV+YygdiQwz8kA8BQ8UfOsc/gNNgwe7jyEqPie7sWALbgUYrAbetgPmrrQxV5
NWChNY04YxsvW3KVa4tOWOFFXAFy9iOcAtsOSlUVrk8TIkez1xbXE3oIP6b43SUePPZS7GVAmTTQ
skiQSeJeR843sTUaxuRBczuWLkimxDnFdV0nru+UMwtSUvP/GWQNx6kWhvJVVXBZr1dENTu11imk
Z1ILZ7iprhErLUNv36uuDYgXC0LrLTNgk+CjcCfkr3nCkIZ9WaqAtyYtgK5icuEAJiI003MDvxQn
5L36CTCa+YEDd24xksOuQs3dzapycPrkz+RgZTcbSgrgcROG6Spg/2fMpoOddH/NoUCFL3e4zbPh
pMUcWphAa7Yqt8z1tLX/NjXTF1DjQFq2Qxe0MCdPKZN2NRDZH67AKPwswwYajcPe5DA4+J84nWPO
TfI48bZLZ0zmf5DuRMo/HcPh9ZpK/PMx1ueLc1mK1cZRA5JMNTO0AnsSLbTb/1POAG42eKevEdnM
5L3socmAPFC5WsUDdyTM68xsuGmsxlvkhY2ZdaXq64h2lDCkGDCIo2n2R8hlakqw6TATVy6iEz34
fsa971N41D+E6GiZIZK6yxo2FBZjRdr4mzX5hWiJzOY7MsiRqz/GVjxjdxB6k05b6e5isI0Cgsyl
MaPHR7gcNBn6+pbhaSixRfL6PUvQXarHTQaUF8N1SkzLM3RxqyGIs7AQ+ZbHtqSk6WFi6Y/r2ehi
bDMQRwuymXrYRKofioCwjv1aNX1p9ewy0PP69rEdYL+sTnh5XHmE2bAnQ0tm0iAnrOJ+3C9845Si
Perks20M0spBmnAoiA+1ACwGaHdGQpwekFV6zzYiM3ItWwaFlbN8Kk+QjsbOhsMan9XXkdQUhl+S
8exHrHZIrG8Lxg88ZIZVOQo/O+XVGaikUc8YJi9182x9llgSmKS79KXO6lxBennnEuvuOmUHGapg
riKYYNEplJyYHlaRrny0csaKQwSZdGv5r+Yb2ekxqOY+jHracoUE1p9bUDCwRuJrlGN+WCaRimvh
XmigKyGbiSsLyI1Wdt5JsbngOeWCJUvDBxt6F7JFLS/P9EfMSAQVAW0uZQ2NC/Af+r+k3HiPnnHI
SMJX8+pTxjqN4rRjj+4mZyhoEY1is9nijVCTCRLNGLYKzQ6ZbNYykhTA4bcr11maOHn/04VADVoe
8W7KTVOADwzMQI9yvlsqdYyj/C5d8A/0p1riaNyUpBxw9FGe36VKYJCCHNV/GA8muHedr5eqdr7I
Ju2/GQ87ZEFIq2QIo0bARECVjlY3hY/ZGUAqh2GyPO5SZi21ZjoBkP9vFOECUgOV9LmApL5EGmrM
0Mvwdq6u7zXG6lttKEgVJVBe8Dft/WNvLxqkLR6c4kGkvPVrhRLhvpdbu0hTUswl9X4gfcsWH0Xg
q0ZG2NSd/JAN4S3/+K+y8yfIEqgfK0nU9uxJP+oYZnqtuWKODiVYGHRiT58w+frlDyc2/2y8DCos
6B3fwIb6miKzqjDOhvO/AQnFpzLwLRT3FhXrRDK9+JwI852nUms0Gc8wLDXNCiXMw9jENWFc6tDe
1W3wwvbP6fk0Xmx4tA2osHPmPPcmncOtVvw5W7WYpt/ZrWlXKFYtaQ8nqpV2RaVWmArP8L/jcMKY
HQpJliSwh4en/9ZJ6LBFiaQ1iWOI0PeOFkd5aTRRKk7QIinJgwfzmkEqQ6OA9t/IASPaLftimOU8
0414SDvmVppamLZyjGFTSBtojMfUP4TUs3Isrfi0tBYTRoXIQienEBNMYiN199F0SqeG0L+ge0bf
W6sWpyba3foUXljFWpKkO60F2zA6emDrt7i3C8HVLIpBIMBWm8FusJpY75AMUckVPxrdTO7tc3E8
DsRMy77qgYSwc/bOkoXdIT8muB9htMTUioIqInqWwrbIgSEk+eHuc2ig8hKYBbvLUNw8jGyJbXMj
oYhXgxyVymPRyJZ9nWUFHpUQFvwe8WUK+0z55jOutot7ntKTvJPWB7aVrsbZcmcwgfIaaHFgSg1/
rDxOeSlOtycqKv4BgkOsGNlLaEArKAKWw6hVQmTYZdvAR+FVT/Cc6eO68gOa6Hq0MGVatuOEWNoK
37C9Fuu3Td3aIEocZnX29fRjSyujnWYiuJPzARGboc8ZqB5Sk22jJij0C45YWnTb+YakyTSVAsE3
Eq7ipz/vHTTOtZx5WjO/O4M11ICQ2IbM07Rc87UkKV/HW21N5CMV2G/KntVcMTd+UoQ/KrjyuS1q
QnnYPoQT+J+91p9lv9LELezlbaG/IfoImXulPnC0iEAtZ1883zzp+3xx3qXoua88lXxn4ziXZvgR
5fw/qxvMEE/N05Ttd4VZsuaHQVMKVXGvpgiur4WNunyw/MW3ItwesQlm/7rwjSF0nHsPjcSHPWPT
f6ymj7R6bNXAXK5Qp6PNAe3UVjy6/aBCOb0XXyjPt7p/MT/l4YselAU7Of3fZdEH7eXWCU6yEP7L
DklV1JHA7cD6dcRPDKRy9UBrOxgtnff4Bidq1UEJ1k0ZwMGn5YU87Sc4ZWimAmYAQEiwq48/SYpZ
wc5bTXnQetf2sPp0UG5p3Kwri4thtTyeGrCtM6TNe4DkEu/ru3mLMoPFnNDEms61lwozQFbG8be9
ffkyjQ5jktiuWTwRYVHQ9EVff6nSm2knLPJAPw90Dib+3Ub5OVBsT/JWOHNg9DiX5rJxaFG6dIdS
c60WIgnbRk2lAn/FyoUZQjWgVcKm460mrE9SrwU/XvCA/Ys9R0HWO3beYy80VCx7KmOtA2FlwOwy
VjADuXdtU+Vml1rO6dXQFiMJgzw18dKOvqyylU9erNyKfXR1nTkQoRVfOAbBmqEh/QW9E+jYqMOm
dMwHjLWfeXzzNO/s9r4cE3pWD66HUjFZW3tpiq/hTwD2rhih+ffWGC+d1VuFmjKNTrrbhKKTAijB
lBAyohgnlBGtNymHoNwgMsG2dlrDC/p2h5gzh69i0sYqehI5r9TMPAFwHQ1SGEmjjws6A1lL6H1J
tg6em8hrJ4sER84jJi4hI5h1LMGC9uyhm9SIzBq/IuJXCESTJFcHbVOcpTR8LC3FI2QNlCbhXD7C
C28nK0OXHfjpwLqSiUx+x9nQ0YplSAwsBd+d8RehYNQoFW/TGynR2qbt/BTgD1YbxLov5JM/6Oap
n4DqOtgRnUwu1GYtf+BXZLeMYAw4XE/bQ2DbHZGzbBkqlDouNvQwkGhhWF4hwYdJgZGF7jdbzFjd
VuWqA0FzizT3ZWP36eEPxoWqWr3xH4fbBybtT5s19rHlmZ1kN6q12R80/QnciSXuiPE+3pFKpBzR
9m4N5Jktkds74VIXNGQ1kbiJo9q0kvfnkcxfYVYA/stR0l1F3bpvY3HOFG1kiLyugywbGHtGWoC4
aMFklSc9z3oZRZIA/j8sjmQ288kPRo+5q89GenjBOBWiPTfiPNqE9FuX2E+FDTje4nVBMPeQHiwb
u9cXnF5/0DQCU+8XYG+6OtGVBNNJKbJWDl5R4o7JQJFbL2XlTRHRFgbc+fyzZUVK8XcIbfXvmqmw
9a9kseFUj7FpO5R3hMVZBwNAKGOAK6pyiyuOsDYF4Ls67C91ial6usXb7ThBCfBmujvWnakdB7Zu
9Wm6YyZTx3H71mQEFKKgk4Y9qm/h+DkS5LdTe7poAdewDIl1epvH51qo5X7rKRiXDEvulV+U3f7W
VhhMT0jbaBpNcKleBjEuFqLkkWA4UiUlXKNlaKrOTwpeWpuBkz9M7imI7FMfdWuuYWO356ioA+Fg
Vu1d9iTMedbE2TrD2emida7gP8ijJA+o+WApIpkgFjD/btC1+vptN5gWvmpL0eSJWpH264RAD54O
HjMde6LepRlzd1OWTsNqQlgwV3PRBTeO3TFKEPouPUWdW1AFuUFX67jZHnh0hz9eo5YiAOpYzc54
/q/lxZJdfUVJAnWbnB4VkxIr4MVijkzN00l1oiEdrrBFAFIf2g8KOVacZUpgjGxTzx7mkXp6pLAc
j8jDdoICkZDDdRDCaLUr9Vm2hs+w4YeaUfpPRJkOTvfs8F9/ETIAefzHRmGastyW9zFOatpI8g9/
mMZBytbTp2ld4O8Oz2MU5D6geVyVgfTVxdzslg41TehhvmeXCJg24eq+n+waulA1aNve+6zYkK4w
2q/Dt3wWpGoI3Jp8IoCxAn+MyjdD6L/461XA3l+0vuyMDGFnuo3hZ9HsgzHGVbYIkJqd/4Usd/iJ
rsNcmcO+mS+BdcRFR6gpUvGumTCWHSx29bYkDPU3GAPIe7+3Wr0PbAv/CJ9hQzwZcnrkXeaWO8lA
Gd5GfvvYSIixcv6zeDUpv7MVp58lbAhFl0Wd5BUrSrvoSdi8QgVkGmq7TvlSqdQxbECr3nhPkuYC
hf4AFopUQp2g3/YaJ6QbWsCro2Gt3CHJ4+DUUv1Veo0K4V/RRsNrv7iQ24+zJS589/yS07B5XMXT
ha9tINun0shraxHoS4n7ADAuyDjrWzGrz9ve7aR+xg77FKYtjmzeR6GMNjkmPEUZ5fx9wzKhUYv+
qI3q73t/TngOeYNes4TsXyu8LlfzJjbZOH1Ahpw/cqnQtKvhf7c6qcThRylw+OusHy68wKaZ4q2n
vSFDeiU7ZD0dDAZL62djpq8COymFzI+ybYSV2OCQDflYhzoAt9Eokp07Nu7ULUDk/vcnqvZBIpaX
E+k9Jv55tenpEGvPxLyGCe3LFfY23nxUBxpmO4WdPBc+yCkT9PUOMKZD45T1QdEQ6b9J7xOQ5E1o
/8ypPUZlOss1VTroh2yfyYAq5BT8a4P8LgonwPyh9vwY54njlzwSPbzvXiCzDWRY1zWGaSjWxLVn
vXI1vWhMLvsk1kF1XpSSUQvurGOgPbO4QmmR82JJO18+XaKU68dbeBnQsehpbPEBGZ9dBAfQ2owr
Lmsa393Jki0DrbxxApV5nENqzphii7xNwELIa7fxj/Z01Oiisqe56seuu9MBgq8HS5Q76Eau08w1
5HtDdMSPL8ZHSwhAhBJIbtYj//6HEv5T0lhm6TDxNJd2ovPRZoRjqwtwCvMZTogIAjsnnnpa9H7G
y3cCZ4VqlGHJPOzchDzFeu9iQtkIonPYHvz8JP2WlGkD+e6xYty8wlRZbF/if6djhQ7l0/gjZYbY
wgeUtnXa85v0eherzjUB8mm1+UywCM64pOw8m20HUVVRTfFC6oDkHjXLWKoC64nMwbOF21qrRFEs
DluYBOzR1bHJsgmYnCB6zwWaZHVpqBuF2pZHrXXcG/cSFV07rJfbanQ8f/z80H/0j93I88aRj6nF
b3iPtvklURKESImoVP5qxiCPHVP08ZTfNyvmPlrKPvjIzdjBOJlwQqUe2mknyU2PHwg9EV10lu4G
3oWvYRDElMtHsZnr+UVZlTn7rep+8phJIPSMX3h775Ij8XUvFDA1UpQNtcWCy5ZwPIpyjE+B34Ns
YterW1xML7DCX5FQFZqlB96kscuNaIoTWY/37xnZX5Rr+T2DQTKYZQThe/2Mz73EmUuqWXNzefD2
yHUmd/at3QMzN5vfoMmvHSitp+yU3VS2pFDF/WvHRhriZe4nWTFbsqpCLcR5fwdAjCctJc6uUsJR
dMwOkg/TDH9cwCK3JLOgIwM65Z51k3GoRyyppjlhT2wCY38Skw68qy5MxLywyUT9w/3k6SoW08FX
f7t12V7VklUEph7nbqRfL2NLYh/zIo4fXo4kr5qcnUQA3XfiJ31jEIkzyvg6hDr0ldILiENcIvRD
7o7kEJtoWNYDluiPSmTd67wS89p9rSiOhIpWl21b6m2kv05DJuWVOg/cn3lNvm48UcgtwqRdgl3l
cwgBmX6ICVPhRl/gM2+ZmWN96bQE+DuwpbuvSJUsIEyJluacR9iaRllqKUMXnWmNTqxB2L3Es9CJ
XtubydhEKYCDRMu9n8CnCn5sbMC2bMgy5UgcWnEGhrJEabJteTGj5RbPrDNu0bfn7aYrJH4sUI28
vU6A3Bek/bocEIwg3mECSzxjcv/ySpmhnlg0tcUInWUNtX4KDbHY8QFvY3UsxPxetsvRGwJrONV2
E2ZhAxnLyB7/EhpEUe0LqcxLdfa3ATekavTwJxnGYf77wWLD0QxoH+WpCCmRt4+zFuzZAw4xw8xN
dNOZRMJYkOCoI4bevGzx78heqwtcLT/LRFmCY6Mgm3x4BkaAjxUKw62tXg1l1owqMRebcUnm84Eh
bha3YtPjtQnwpKeTRyvPakW/xsMW8sHVUfVAAzKqOTOr2gEi6spV3+1CGZFZNXN6yxksEPcv2zEP
B8E/E5f6EVGcnJ56DM2FlUj4vxCLEbWKw+L7UYoy9DdziTxQWWm6qKLOJBHze07o6YFJag==
`protect end_protected
