`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MkwPv2wOZ9UXSr6u+NwdPbGxCffbA4pIiDeEjWWtF5fSpp6QZrXVsRqY6/NthUO/iZhcg46Rng19
qr4EysKP9w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jkSsmmUjSHEl/UhliH0rvSFNUonl7+x7733ytFOuwlKURjmkykqB6qf2F7nMvtb2I9l0nU9ut2YU
cJxt5qLTqiXf9VyYxKz6/WrImwAMniNkvBxb1jwpwBHcQaDeIcM7hz6woct71S5cPmsHU7DZ6fP5
l8R24zuCM6DosMl+/pc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3IXM5jSYeJWDSwx3PtQCBsDOv0c4c85w0tTiWFhpMp2htZIc63xXBP3WHabH1idhfVk+AmLhLCCF
flk66KtXnWwancYkYRuKWhrNHE+hCXX3+yVnMikTwfCx5CoC+C0WrdQsY53xbzoT6frMUP3nm8XI
F5JA3ZBCYCBLhrMjMxMYINCvoFrKaGoI5a8WSwSz1aVrXbf5iwCkwCrAE102qDXekNE8XBzsZQ9G
0x1cgraYom8axqPWaBsCA5cXPSzZToRt33VJxYK+5z1/kNhENmL4QAZFgc89kv/o3jBqyS21ffdR
e6esrHmUB+q4sKVICo84OUxfDDQkqSTj7jmHnQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0PU+sr30a8hrcJpv59TYeaVTcNUQhQcnGCuN+hh+/hlHyv8oqEL3DMo7wVT9U5mfzj//R+m9kqI6
B7NrYkOeA4t+XOXVWtyd87kFld6jktBzJ6JAygrUW2CyeCaoSoTT8mlnwkEqWZaZC/ET+/Popfsd
jcan7kVOB0AkTIzocE4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AuWqOtCw5UtGBKfYQtcOKMNqDt30g47OeqIyTs1u6eSGPppqG+SD4jD4zwOZK9jFP3n2iXznzGWS
DpOEIERFEOJFnenOFWW49/p6z/BnZ3B2klKGIhVv9oxVEwFZqhS2q/kp253QoXS02xIHKQVFA3Wv
RfMFtIJfap/jckAImS+9Q1C5iWy84qUfsueBR5rNz1tWhJNnMkR7DhCtA2M5/bRL+BzXs7HdGXYM
lcIqqiaoj+XTwD12OrMbMI7egGkKGo6HAbdXNdtvuvv9D7vAyET3q2pRdlBKYedAVYC3Rszfkzr1
ZVruUdLdC9IQbKWHNKaP3Wk/zt6i7/oG2Gq74w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10432)
`protect data_block
VtovPVrg45oeEARG9dWm5YXzIilmoBaEhO4m8N+7lL0C8yTv8hb0VRdn+e2BGldDVHE224AXLIuR
aIC6cEuUkyY8CjVQ8mzYBjNpWBBM9PRQ2KJOSiCATbvLizrImgmmFR2+8lFQVu6Xub3kKmfGt8j3
asw+L4dn5Gvdw34VJZ4/eWeyJua60cjj6T6/DnvF21cHFpKZjR1veqgbC+P2d+RwTXWXMlDXfS+C
wqzleQn+jFTbRyukWt7tKsGuOYJUFh0n0LnZllFX6K+DqnEegf2K+k7iU8QMcZmMSWseCgRyfpIg
OfvvPTh/WVklPj4qm8fcFkgEaFpbCLoofbOn8ALKW1dhH2TrUGh66OHusAePcOiAUU3lpIZppMxU
POwevubGMPnX0BXV3YHxn8idgXMs+8Uj66I7zA0rQLEK3LpF9Hd5kGqYItlpGPXq46KugL/EYtqL
SqSUR+CL8mezTqeCIsZX442/jTVtZ4BG5qt8kmprJLvsj+AN/FjfKiQRwRkDuaAhK7l/G7+UvVjJ
QRRDGB+aaHu32bvrf02PR7bDbFnybdH7RdL7Q6sfGhMQNzqXqvbuk8WxIHp3nsvTnAOj0NFTBov3
npBrtl6P44vIAjb9nM6aQmtC3qsloaEk6pLwtgCTJBjqwRps/S80OlRb38joE5iPXqnFJlWkDtlf
ABs8VJgA1ld6Utv9ScdowDf77wQtTzT70PFRC4gaTuscrzLADaF4D9fwhj5mpgV//3nDQFjbFrzs
ctwVriGaO1LiW7Xlv0F0UIqcfNPV1KURiN1XYBW3/O3jJvtIk24Oa4ZjTwkgXqDVubd3lTAxhSyj
p2czZLajbWL6pEITo4dQY/qRfjN4DRv65dyWBafLcrXUxoRp7GROdoT4n0wYalXdmX2whnQvdio8
55cJX+WIjdB9FShEPlnrcWrhPCVpSzZxJpo4YPHsyYpOS0PSHvGKGAAoEaPjj6Qfx/lEwhf9c2H2
0kHKJpooo1WOp716tg7OvMe0Qx09mt1MEK0qf9w+yk1M0O43F2qqWU6P76UYNU/zk+vABw5PHZkl
4WdaHPf/npXX2mTZe8V8Nn2/upTc27749KXLk7hEuDlJU+eTB6bnYtTVBRSQ4RqXrBOROkvkZaFe
s0ZUq90B7TgoX12znTCigP0UyPCq03Qoo/jtJUVgozLP0O5M/O2fGHHMPO5m2JjAWOFjv6oz0VoH
fL4rCaq27e+Qc+eKGOwZo1BZDRdjnF1gAH4Gwp2GtzFnU6p4P/HtZGWYXF/5rDQ0QEv2coQgf1+3
PPsAjGLkJ50orWrFuy9VKy2aUMy7s6LTMvTG/hwFgmWhgLlYTP0jKA2npqdKk9op3dBxirBa2Y+V
V0ZOzi7fPL3AixFVP6eu/HAJFcXzhhoX9bZ8GMcxPtqf8W65luIRztDrpMCwvJyuoVF4/CAu6OCg
jV6bEVybTSgavr6RNHkOnWGRUkK4dAwuep2YQjaU2QPJkl1IqO23v0KW9pZxnj6CNXARSrpXE7ux
x3XBO0kfoUnf5Ic0y46HW8Wb8Kp8HInEn/EJkhfPneAA8AFpZBXot/n0CnRls/w+Ojp538iLFRsF
u9FhnqUu5Y2gTViOfipe2x+dSTf+Q6cSf7yDLDWB7edOP3e19+rC6ny/hgRg4aVkPg/pQr3ULVtT
gY8UOyW7NuDWUtrnObNdg2GfmAeuKoos4EtpERnKKQ0s6hv3bbLzg/aEByS690C0U9E0kVdm+KT+
pq2tWj2JImn8YHNgegbRiqTFmjNfermeGzKpFgZJrQ1k3M/5lhVjG9vkyWWGDzuLX34wSkV09Diy
fEVczQnxbo4MIqGHOsdSnjEEy1KYHeHW15FQLdXq67GNdNEBj4DpJFo4XjOklMgFWjG7sYeX3fXP
KHIzLzL/hQ+wQIoXhFb3vJUXbnG2alZgZGyC9dvlU4Z3x/fsibfV8x45/Itgbnd++JDIQn6HXsnG
UjEWWbYg+VOmpJbV+Fqj0HXKVNS1WmmMB5Xq6WMIowxy1/2pN6ZEF4vKiWV0FYUaJhwvuglzk10T
cq00EErcju5wv0zZd2LBNOs2Xt11Xa20R9scySA9EoW4XlwiUpWVXbQFcn/8aX0w4lh+2qL5nY0F
OAkMqcQnjtIU6SgTPUQrc/fOfPH/zM8EcGIoQwb9NiAfOKcmHqX7XECVAEIvqYbVMzJ+3O74YEH3
LYMAP6YSrQaesOY8aZqBLYlD2hz/r81eQO5HbeqEo34jLynneYGPyyNTv4rJx7dK3EcCMKMZRRRv
bm01xpEA7Ia+OPQoB7k0ibMAPrhyBedrIit/8Dk28sM1HS0YNzZf6op9pp4X1Pfgi8td/ELeISYC
CDcMTt5Z9que+s+8R3pcfWZVhEyLwSdMUad9QUT4N+Y2NLgC1+r1Q9KTfBCmFTNbSnpzJpELQkQE
mcopI1yJexOLEFeBL5ZVLxlI60aF2qFNP78WQGdYD7Zt9DoQ94HiBngt0epdDMuF4T5CXyWb3fmC
hKNcp0NZIB/g2a5xRE6hUEOtVSo6aji3UBO56SIzfimmDsH2xfm+0jM2KeqU53rLi+J7eGbjBRdr
Cp+p8UNSHGZv9CrQXjftKxDISEENKsCKG0G7B1ZKw96alzCAm8wsLQejRNZUzvdAKZAYuweWUm/B
Ken0EaeNKkQjyYZR5qL83ekE54EFKcayA7XPggK+6e5vK76t2MmCG7DwtZAjwUpvJejDNc7u3CwH
HNTBAzFN4725NzKM8xKqcwfcK5prkpPdNQEiVOMf9+QPm/kZJHkX7qNHi8IAfHP2QAL0ZMIg9urd
1w8j+0/D19dnkogkN8sjLkCP6TGnhhMePzLWAwmeesIt4pVtiHeXpDo71DOPCGyXr62RHwwJua4Y
oapDxqfqhRYvVQn//jeAHRLjHMem78E7KWgZ0rCrS23F5fPytNblgv0KQVZ3Bk7WyzEN94l7nD0O
n8RKPW853rXkM1ZnggBdBjYcN4QnpVVC2n/2D5IOoaPkOoU+sq9RSVtCMwh5C/C1mLjonADLpIdX
hE1S19AQWKc5ESjo53v/jR3vstePeUCuJW6CtPEwrwhvH90a3vryl7TulBdohmGqL28oq+8Kp3WS
HjlQXhITBm/Xl+uA0ZCfwWKsuxNr24rOIBPrqvKEaZ4FsP6HwWJi32zSvACLGMbWjV3aGL6Cx3YE
Sm5BrL+s3Su/lfU9b3gXGAMBTLMzxJJVauqmCqkhu65FQW/A92gmRV7SjR6XHLjbwFHn3ybRSdyo
i/+e43pJf4JGfwsABjkxNuwrjuonr/FEk/r2XS9uf/BmsooiW1x2Kqp3scVceY/SFnRLbs7l7uEB
1XrV9eIv7Gypw8K7uIB5S5YYmI43bDf4vi20QcRRsjUGUaRHqRkj4AL1P9zGawo9Oh5Az7HkQCNw
OruuhG2PRdRm3Vs4xpfHgezu89PYECcklmkff9SN5HBK4k/l+5qp6bgSyYpLFyxmEo92CvoLXGPD
bcAFE6F27b1XTqle4GDh0GbspUnL39Ez7Pdrnf2nQwbrXYx81GEymxb3pPEwHo+XnHxsI7v+D1lc
09kQVzSJBE75ZmM8sli3EC6EOuLaWzhppmcpMgHZN0cU+m5vu2EoIlEQPSHCCccZGfnLwOhe2kid
HbB0kcOl9mnPuyr2BN8bcUgQSX0ft21Vg9oh3BonN/vMyUAkD+ZuPGVqkMKmv0pm3Nx2phFmkHiB
2w3l9ckp1Cmnt2rITKKRZiJOBgpQ4k8nWx5ZCKwJi0JlxFTIqI4enDi31+f2CJNN0kinjVB1sjjM
6ODwE583yXvkxVkhZLLxJSfmeGKMqjJe5SoL5CIorpdVUZhQdfO0ObEFcg8Zsso6ARoTpn+s/lMo
+WI9k35QG0cuEwcNBQDGVyasg96smSrSbqAawhyWxmRjZSyA9JcUmMoPt3AvEJKoyQUjhfL1kgCK
E4VBrEOog6z5BSsbVle8ksLK6jF/Yv/ZGwYPhagbI41AuaY2Cwg5ArxHVyRwGfAgb3NZKV0KFI31
eXgy16TAx3on6fkM2ytYDH4BNCw6w/cMMlEqUFQm7JtD4enJXXFp43rzr18OQMFNZSEV8/RS7Xdj
5kDKnccFyFP13H6tw4HRHgIgebO7cVc25C/ST+BqkrAv36gxMLgd8qX/tajmlVV2mVNcFiGFMPxJ
AEEVh5XMTx76VkgOh4ReHiut7IgZvy+yqIaKnfaE3Im4N5CqNuk5U39lfRkbmwPryVeMd8OIoEqQ
H4CWHR5i8JqWD9EFWMXPFXC3Ntg7ZzH/c+31MG271MqKs55F7/3FDavEjQT9BO+oBV++AnEpSfRx
HG/3KyHQ+PD4Zl3aO5JuV+ec/ggGmiH+8X+Ub60pxtOS3A7uEYHqj9k5t7aG25i55MH5MPrXEDRi
Hsun+pir0y90qftRZgu2Inz5bbtQUCHMdAysssxRqljK9KlHAOAdHvYxkVwElhKzi1FlNB8ymoBU
GRX7Wgyc+CPp4YAqyNpUyPAYW2Ct04rSbY9owxMrCVIeOjL7y81Zbd+vgYl1hOj1JH0/Sew8g7sp
JFjSgIrPgoiOvQ53EIghIvCmMBl35jw3VV0GQQrt7B3kKgfK7u4m+pTLlWhPZ1qAKER7QfjlXuBI
TgOwDoXhGzzKgmgzk84Jl8mLcwzbnZSWxkIJYvzG6tjCgqrASCn3eXtl1CnhP/avTXv4wtiZATdz
/rqdOQ+TWthJ5nztGhjbSXuwp96v3L/WOXMVTm88LsLSJKszIb+wKCmI+Kh6I+zo9jxCn9AHnRgv
f22hp8OjnPjyQsS5p9K7yHpRz5SwJbEJkXVbrQMv+/JqSxO1nDyZPUdK0rR1bQrWnOFCLTpoTenu
Dbizn650XWEepw+xdmWWpfLAQAR4BNncXOSYgkOtjAnOu39X8djX8Uf2c03Qi6S+LxiDuMUE4mvG
4c+Gn+N7bL5aLRJ/h6b5m6ao5P3R6SIgZD7KykknfsHhBzFSv8s0cDu1iE/hp+D4TRSJEJWaYKAv
dMi5/5zbbWiP+HCZlHFI4VdWBX55e5v2+aHq02+EM5YrUfG4wjMzCa4Z6xSXD2nhdpaI36YXf8fn
PWukG1RLDBzf9IykzziSpSTmAbiKOw7MP4tJNMjepMW/1xXpb3MHHaPowp5Vh2ENyD8y+7WEy3ox
z0Qtze51ZDp+xe3z3msjsB8JnaMYwDgvR1TSbdCHXajABOk5HIvazkQYUTON6B8P4VOrDn8ANQLi
6YEZLdxPZ2MLmpE/3FrklQ1G+KTa5ygP1F1CcgnaZN/o4nLqaI4qpGN030ysWSEoRg/KNNpAQoqS
T6nkjgqoZrPSWu1pn1RXY71+SM10IHDLM4N7QrbPk2Eu2STdf9wSJxVPjtA/s9bmYujOhGsy4vmu
/POzMxgp4dc9qTcuPQnGnOWr55jr2+YnaujpDZw6U4NDnx1CCg6PNtlYlp3rL2PEu2BwgQWCffAu
k1/3EmrLlIijdeNcWLoGhUXmsFlq+oxtOGKhCiqGfKtqZuB4PFX5QGwSPbWkc08PY201WVdQuA5q
vdRcSvWqCNNQ8j5i9yw2cpCx1A/mgpfBfXSz8Z3pA1zwj7JOB5rBlzUtH5/GgWCg4e4zEb9R1j6M
LYK6Bx1u76C5vHPmLaPkokNsWSyYCTUATzKH9NZwvae5ZY5ttfYpVpfTwEYo5/loSFE2vhpIUsW7
ycsl7ylJeHLqwZPhkgWtB12xrTV0M9TVuacdwogq09eQ7mHBICSMOenyOgArxvuGGEJ1gaump7oY
iPHLTiSDbORuHvPkHE6EVKch1lHJ1aR9ch6ba6OXssPUU0GyS4dmv6SEjK472futcOokpoMQguYn
7OXkYtYiP2B3YznxmjNBqyvObesZX5FdaD6W6CL2Bjx0818Gqht3keiZapJNAxGsR//vGTX+DjbY
Ah8Kze+HaY67KMQMDc756FvOrWbmBjcy0E2VqgwOozSj3qNNEnAGUUh21p1I1W4sR65e3++R76ZO
q3M53ALsiIhZXGjuzrvWa4S7kJkYrEsryIjW+3o4feQ7ZuFfux+cTUnKwcHSFTxzOlLFiDelLeua
VQjd87GDPdLR4phM+5dq5AHFSKoRyAe0/e1QDu4iRQDmmajY07xOV31zG8S6k52rjtV1HB9rym5Y
Wm8jEL+ar+An0yquNKKPjjxU4310Uid463GTgN0IB32c9COU4LxWsxvtasPa1uNT/5haFOMCDPzv
au+eCIS1OWcY1CU2A9Tiz/FNsI4xXSHk30M5OojMUSsuD4ybyR/LpbDyAUAO17vTmwnsNH6bDo6H
hkJilJlrUMigyoyaWGwsMVymRPTYDJV6nfFHzLng9pXT+BlfJ+LZUyg4IkwtsuU/Hshn2Iml6Im4
Dfv48PdhdNcBHUX4Ql9mpS3zFeDeaEKlWUkm4fBcjso3409X61ZiDY+ItCgSQkvYPaO6UllPBOiY
nJMFj9bzz8Z9ILddmTWtMVR33bYFAzKWALCxgUQBft60URQ4OhVyzQ6/inffmySPDvhDjS4FaBvX
lMSONNPd8hPSyH/osUvV7jFkrTM22ZXwomRwBQyVR58XunAPyV70E0WGxQmI9GsZdGfqQqZ65Wfx
Lgzcdgzoqlfv6asMnUmFJpprP98kXy6J06vKIenUKR+aPuzPFMWszIjRHSAzxf6xI02pzamljyzt
FYK7DZR59K6LFR94B7FooAQCuk4vJQ0k2G0lcbd1RgfMtfTR/17o8VnrbjquktHfGlJcFtNm35tH
mzS4sGqYQ8KkuvJYCI/5+uY/R942jzlAPNVl/bgQo3xtbE/JLqD3bzRbk0RyFVap+fCxnklmBcXb
HPf1UtAx8Cgwsftbxnxm9n9jpr2waGml8FljWu5zCd87/oBnFP5DvM1PU61Wc4jEuQhS0AgnCR7d
qywHFdoTPP2GwLf3eu1VcfMe28Xg4Cgcb/p+g0o0eNW8a1ymBvEWsJx1Gk5Iqy2HmaKX3yCF0yNV
dTWRra9OCIjYwONncuUfILnxaNki2fC64IkqcIkJ6EGbIyrPEHyegyNo/duq4rrT2pVIKjmCB1Rw
afzVMH6z6y5SYYd3rq3rX4kP8+IQ509gaavv8mRQp3laQ4tBymkg3GFJwbWSpn9R7w1hxKPDUz6q
v16DmZjiNBQ2LbUOgTfFruU54y2+K29f9RlEpNLs2yUHgBkr5IW9CYmP7iuGqX0cOMtK/Fdu3H2b
sLnMY0yfAw8Z6cqLTeOLGQVaAkKv3nfN8xoT42qb32Gk2jxLs7LCAlLgkooKWVduUiHVpm8ikr2r
GTRm3l8Qq85aN0IQ7CUQc8tTW1YoBqkNQ4SGWpPH2c64H3/FQbwBvZ02cgmpGjgkEXrCmUKVZL3E
QH6RKmMTUKoywMGdeT7qXHs8k1rdnUfuO+vogvzuZIfT/wS/gjZ7Swvsiuzf85H8cXFhduu0p6l/
O3keWyhLRDlrkuPUl9DCk5fQGKC67Qtv24LBVQ6LAN0cDZb/edJd7F/Lw/nQmzecrC2Evy4nZ99e
cDNt2ZvsBrCXE/AiQXK/FsYU1b6TVbKXRdEG31l95j+ObCF6YjFmhbze+qW+1KLKvYjVFvLEPSEm
0+9KrkbO4HlpotQk+mOHAzHMUiHW+J3KRY9Q5KHeJzGh/H+jGlv7NlcKsfBAsEfIkLAqSxvpNpFJ
1Xt+oGqc+BnPVMPZoGpL2XxPqfsMt3OSaYbBw/ffPnPYnzMJXcFiGH2LuCtrveqU73GOK3ZKpp+w
pcCMSo8egBmq4Ve4SpLe0Ew3f/oBdKwDOF6vcr2FOSmw/1qg99XoWc4Yo36NTkjgkbrM6Xbyy4VI
sqZDLATZffkjew0FYkNf9Qf4mQ5AMOILQEttEiI+JTbJc3ByemkonGppUREosbOrXE+5TT78wslS
rWjc1VfInnWJ4pWrFgPohbgiq9reEduO6Ug/V2SjzlZQmuWhrxbFYSfh4VIjWcI3pLFxDkQiOpUw
VDdjnUGkIc8/Lx6zB/vlpzTF5NkREOn//BGtEAEQKBWVz9IyHoIzBXBMjIa08j15CaHWv950Wa/4
SelmZHbS8YhHtGWjWpCgfSy94H3AsKlRV/wpUW6BwNKHSr4xdqjvDtYIQTD9YvGcyqDffL1+gC07
AsX0U0hHi+/qcGic6pVOKV21deFy9qzIMTlrFH6LRr1JIKOmqmhWdJIgNIusIWkwzfVvV3P9iDnH
o1j+cBJ+uLtORdNmGl28RSIFASxv+CgVANal6SFBdvcuiXRKHEah4Ug76MZTNaZp4AGPbLhTX+a9
LIZfiy9XrYTL/BOxxJW68jJNSvj7Z0usfsxXn7/UwPVtUdJOroRL2PnIMCvPiWFPs3NLYj6mnr4u
ud33JohI/j+r0fF/HwCovK6rc8QxZ/HlGhANBuqDwUCbgVjm49KDtxMy1iepPbbmZ1G9p+OASnK3
1InhFX6RrO4WeNPf/wdd/KCR02HO/qjteBtu6+o2PZfmEQ1+J04rJs9t9eWECXyzGnlW3u3bs7NB
BQwVNhjvKbWtiRyCt1OuLp4UMP/y4cXZGW5kQHN22ZxEdKZFsWmgVeVcLvqLAoc4zXC3/wfTuQ8q
PCtMRVx+2jZJGy6mLyDsKMbcs+K2dQ0uQHq3JDdEVsLd0sARicqOICNP/hSDlo3k5TJ2wQd2qFGu
e/iAD3/otv3JFLkHaANfChw4C6SDWr684wz4Pjh1Ajb3Kv45B7mgQ6TYl1LVOekEeiU92SsrLzxJ
+Gw/m0SyZWJoWRvs0ReODz4DjLzavIQxb1v+UlHF08C3ZS7EBzpyt6oUeelXzXKqLFdoWdv04iJD
irZ2dZQ+AC9NoQo0p2S7wm6nnEze4SHpD1gUox10cdYzY+1P0dmR82B1w+k/LJ9cOCfnfXndtM2y
IeiWFItP3MhrpIQU3wvREPFe/5/LmXXHwZxfTblxgCqdTrL/paa8U6iX2TFoxjDz6p+7rE172QT0
1xKrnGKAHbMxLmAw1/CsgOR7tF9xBNmeslIyrNMP63PsjKZWOOeSisnmyu0rbPjCzVDZjmc6NsKc
rZd2cefDtVzoxAq+1fSW4ybbGRVrV7bWO4MNVff7oWcWndc80rANpMoQUvyCUs0XidzyZ5HN1KGG
6J4M9laC2wOrPdkQUN+DERh5SFw4LGmqtMwn16Miss4lqqo0ddwjhF5bijsLk88dq68tPhuCcntV
A+VoP3XRwWHFqoEvqEz/z/01nErVkdV/Cz1doXPQHIilvlxFR3zNGF0DhmWZQ5V8lIyPxmESg2Eb
fqYAbz4wFGSk8txWC+0S/v02kMpG4r2OKPw93+ZF+YCDU5FTCCkx9avHLB+4mS1nbOwIyP7NR0w5
Z5+Bmv3wckniBNGNixyd7o9qFjP0lTn4z0kzWy8zj2XkpF+S0j6hk6KgiaTM87An697QOJ5phQF2
DUva44rD33B+9+HVgbesNt5PkHMN/pQd5MEg7/f7+nlXMG5IQqvbh4Njdr2xsO0jpobQoXU/2hDt
gkliIXZY4YyZdKISv7hRVTDtlVAF3U1JtmHsZhz2nbepUSp/tsGpeiKtcN+kFnh3ajcwmyOT2FV/
zMv8IaE883TIjrPBpVTLAk+ReiIzzeTsjD5EU4kt6OgFA1LmaX+VgjYVsFMNsFpFy696wQHoc0G+
HU7Bnejd+8m9lCj6qN2ShJzaWdMNZmrUx3jI9XKP06P5TaZ4HaLNEYhVc8EA2uFAJGUbrihd5FS0
NYeO61MTQbn1fsJHE6i8gNP196SZSda5ElgUysF9wbGORxT39fCkwv1Yq8xJK1ve2qzEU/w6dO6Z
xPhziENKz40G2lz7eXyM+GDY1R8vfcuLmr5JlUEStjuw11CO60T6RX7DobG0aN2r5ZXl12xOmymq
6UWMAu16OfpzJWK4nO2l8NWM2akHbo6euMyHQwk53yXjyQtcq07VjJTYLP7JsaQ7Op8MWGGeRZRS
uArdLSX1Xw3ZHS2V97LX5r+/KowYFqxQHk9hfYIJrzeMhaPoPZGyqeNMo0ZARIKt/ud/yP/O5jxj
SN6gkGYRZTZDJ3xoR12i35GP1Ecyob42CCzPw75hNCaXy9qUAq7xzBSSwTV2CcHObzeFf9rJotjf
ll+lmFoKhI0+YYLnk5aaTlcgNgs2JaMFTHlEIIPywUNQcQQywvlfp4IYMT12vcMraBygAPrj7zo9
nQj+O0Z/06+W78MuGb0e/bNgTlSxR8nIfxWh+sKY4tUVcN02pzvWPfSrIJxElazT5z3Hl+S9/fJh
IXUK0yeaU5LibZUk6fzUnmGQccv5NkxfiI/nf7HX8kdVzXTD4JxNic6LU/QhzuI0cplvy9R0gpIG
j5JxzdsdVpGvIZxBhYn6QlOJbB1GZiGNE7yOU6heLWZZibs3U3USTKa+GBeCo+phd8QD6g+GKY33
45Y9nBxDNxiUSS4xOIDTVG4Z61Bpwp8tWGWJDJpd70rCJ71O3N8jCmMaBrcGH/7gcyinqRWcMpWc
RLtDjsEvX3t6RkERbVM+J21wdcx5XVa16gTSFSafc6rkn0IXSsfLPpiUJHQ3VVc4oQBfJQxeDuWI
vMoyJ7bwqSH3lvRPlZhp0rvxpR8lro1O/+ly7Y6iCPG5Z70/KdGaV5QJsD3AB76IXRuj4wWdj6gM
wKBXW6i8SSuuK5N2q0Af1VsE6U5zjEK5kXBWaQbAK4ciYk5bJ+CSAnu/APesUkk5RxCZiaRqWVrA
xJYQt7oXshtwaD/n0OsE98iBM1WWomFA/3cRFI81cj2HbmSLYzPwZ7DBi+nWVoe8mnz6vR0mfL2p
GBWwj2lSSEZ7LX0GgMB3gR4h06XrUUwt0jTUkn7sdG2rE3WNP+zhE8uld6ha8Aukag+zqBUToOpf
yqzx+OR0O5WMOC4MlRbZnSh8ZMoy/WvLOX5fE+CYHsir6Vt9h8KxyUbkKZbERhVh6lEkckKiaNR0
hl3mCypp+egDBNa3SC2paDXxODYV6AVO0C9PZVskqSu0jFQg+SbPx8VzS0jraPEIHD9Ji6Dy21uQ
d2rR55T1uly/qmdzE1isO8awmmKASDrgJVsuSMcvyReGL9IlTrZLG7oh+ciKOCSD1PHygkUJAdZo
FFf8FTfq/RnSITatTiYvkiy/PPuN3FBUJDoDcPb7wxS8lChuYf9ALcOZMNMuwRxEZU8yefa4mRDP
pg4Ae3wocpHiA0SmvTo2x2STjaD5EAn3Dn//qwp0M/watjXENuLjlqqwmgFEVSySS6uHL7N5FT1K
YiCamtqjf1Sy3iJhroJLFgeHjucftSUwY38e2wt4XteQvRZG3zY9dvie0k4OnBdnjQuh862Qbvi/
ukF6E7GZsGy+YfowEg2/MstRPUk8CRXubMWpcT5pMFCZwKXlAUpP6aUANmVc/86tu7mHq2Jicpcp
Wo1aEHeDz1Hy9+pt2yGV9KNXgzx60ZY6N5tMs55/xeKuPf59x9B6DibsTUmt5G7nYBBPKts/3Z/s
xQ4a/ohkHDb5ib8Z6L72BWbpUyBQI0oSP10ck8Y3wdZ2lbsGE85ICPTE7ySvF995osh+QUTjuZPQ
t5t7hDD7RHP5XcHWsmQIxqt3d2OohS7N8ItioEunvd1+k6LhUV4O+FnHAVBEOjQuuBtoC35EclCy
Pph9UMPqAWdl6nsd95d7IhIJThUHVa2/om9erZGqNhDv2SOEGDszGL0/R9wVSzb+gHXIv+9H2580
jTFntA/xSWGebY/deGg7o97IkI3azusb9/xkSayRCghinVgql0E/JuEve3KfTAdaeqpbBsJsFcVP
FQdZMH36g7oiJt0mjyoiRv7XmxcPWHsz+fUvTFHPDfwvmx5JZkk8WorZcLFpGCFHn9PZg5Uh7zBA
byRPX5uGuoPUBeiX3Ntl/z1GrjBgo5ZKOehN5gu/VZz0pofL0ezwoHzkbO069D3k8gWaMlwFf40W
1pHMCwDHacCMPviomS0D86HLhoI8XtNoZ7Apvhk3WvbOkL3B+CnKZsin8EoAFigV7v22DWpmZ9qr
RKTGAC/sgCj7IRlXR1mgwlZxDDkn+m6dRSgh+wCfaI9v5FUFk4k09dnv6dh3XRhQWpD/ZKUJuoxg
PgndPS+ggCGjY5UykQN6EH5Ys7kXzH/V85kRvMAqzEyMyt5OEaMysHZBd+DLY839q7csGkk7yiaw
quFgQEwPK8sK6+qklpBFTjX4T0AYLa0VPTB2A3ZwF3J9arvir08yDgXHED9DNNVdAD7V2OCKIJQS
DGorkIQOqTtjc+kxX2dqTuTRcztry5WRvYIfLcrNP3ah87K+iwbzF4cE6/NrHkEYsm1QY3qFLP3Z
DumbOwLXc+ZoNursrzcJV9R3XJ3o1hEJI+SVbWtvoao9I1mJRk7KM2I1KYoY37ZvhrNSg30rDq+b
2R0WMniC0lF74s93606pPsm4v1xvG7QF31FboaUkoOA+MfsNHGNqgsGw1ac1em8Zvhq9D6m2IBnb
uUtQfJIhuPankq2yg/b3P/pOSwiG7K3RscCDXlPddSXl9lJcCNoXH9pUsivXa+t1s7T0fVLaYMrN
TFybCj6UbhL+jJJwxlBw36PFBR0ecl5ngtE6zA2Rbdzb+CERrBFQQDQUkuDcLOghTB9WPpu9NFDv
dPSjgEv2nUfFwA6vF2eCFqjvwN8I02sZXYLBBHWHbdYzJgBxSnQBn2aTa2HW4VYXwdpU1+pGgqSp
4H/CbImCiVb7959HWinB8+gw7zwO4B8Lrm+i1NeLyMLqCdQMEh59tjZzLftaiRW9c5mSmZjNU9Pi
RGOBboQdHiXBRlRetO+yHJFDkIra6fyQsFiDAa4M0jAyF2PiOxdnWqCLy2E+IkUKdALiYSeXBuad
055IvMKDzA6bG+08X6xCcgKAAKkkcO+ZZZ4IRntIXupCCiGkQCF01OK5GHrjPb7IJ/hPexZd5P8Y
oJ2Z3fgcUzkLRBUMTfMkpHxXPnNBd704VBKjj3bEmFCEGC1ngdH81DnGuRF4pqi//2X1pm5FXuIy
FCQLI2xcH+orjxrz7tTyGimeRtBSH4rB81YjkKvMJFu6Ixwp6QBDVadmOZlmDtMSvDsszZJAFMNW
UQEMqdHTR0SCNb97EttVFWOyiQlGIELkTAI8c/WmBUyNU+pO0PyRDXgVHjrgKJkh/4sAIKlo2Tms
/4oW4c5Br3ZK8OakcFPxhlVs+9IE8E3EFRp5uLYHAab0sdBGTlX5dELvI7GhGdoMVP4ZTZALjytn
HAc0tULy+12TuFbkgEflVmZyWZuCyED3zM8xsbwK2vVmec7i25bdZltNA1cZ4qFwcylnUh3GWs+M
ujeQGB+bv2bhh09c7YgttC+VKPzowe2O5eAe7Emc4gZUEluXDcpX5VVy451pz+vwWizeoH6wFsfO
RJ2d4Haj1i+tAXmqOvcl1Y5MKpjb+nDmRX67ZM9s214KglJREOLKafxKh8WM9eWjRr6uirD+ydb0
AJOIFxdl5I87PlBl/kgLhnYO1IKevqL/PHWvHBjEEVUQvNag5xKq8P+0eslMFtdoF9JXHxjBrh3o
t/xHn579cd4zPa3ndOjf9TpwnLPurlF7R2+feDwhxT7kHNCMiUM7Aqh2Tw5MvJrkoW+6JnTOfpLV
ue6km0hnV4hJtVctW0WboYiTkJmQl3mBw+KnttS8zUBvV8xv68MFQKpsBaGrmVuU42HVdGuVY6Hg
xk1OR9PDpWakokMyiXMQXXEWINr1Sbv3wfZ2DuyDCcCg1P3FTWUvkjaF1l0R77NpJCcv5ZAiy4EH
61wHolVLYVXVtIxDALdyv50fYDRuyH2Bee1klfPTV7wdloddCQdtqDrK8TnH54acBGLlNU6rECCl
sJhrgWqfC3G0PBGpdXMzHH5nj4LXIOV5x3TWmTQtG9Miw8kr7PqQGBq5hUO5ZRcBA29/0Asfbq0h
5Q==
`protect end_protected
