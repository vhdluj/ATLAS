`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hrt1yFpMpSI67+kaY+BRT17Qdx0DcSEyu3f5hg4VR2hFLm+DdNaCwSt1Gf4oyt6pixTOp4cHWgY3
rvQR4w6EPA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nBiz8eA9B7p0ZfKZTkGApaNvbYyqluwvDYpd7yCXFPVRCDVdFkOk6MdW37MfuJQ2v/ClZikX3V7Z
OLiVgkmnmVAfGJEF8S2+oQFx37hwTzd2sKYiTATeTaU4a+LPNIUfyUkV2GmHEduiLbEBw/rwagX+
P9CZkI/n2BWWiXi8QvY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LmSsyA2TWcZhv8y0rGgiW8QtwKX6HvWmHzqc9Rz0wj+C3rL/OdmS2WtmGm7BhYBMlBlS1NXNAfFP
0E0DKLspi9Cv1zCaj7GDaySGIXRkhevMGxDzovXC/vxK6/gAtcEkfh2A9gegdc7DlrRaZmzBkIQH
xebbITmwEaOg+cdOkZi631xRro86KI1sPeztSc+kMUXruAoyWSsoJuXFQpUu4FYj6V/cqCOHklnF
/+jUI74GDCoLwENa8xfROZrxd6WNU0wwonwjLDLPfGMTI0ZpbSspZKwVzld4/X9GDo/vWuB8S6X0
MTocY8xefNqzi3BmJzWcrjIj1cuFHtbxMUKZZg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wHD3RAsc1ilFgWB6O4vWDWd1+MszNZ6TYmec2N5r1mHQTXyzp+fu+zyZ1uFQ29+Ji6PuiJGLeDXh
4AmsoIyhYP6R57UO4WHpUgCr1256Df1j4USkT5opDtZ3J0AUvf196Fj0bq16yFjYxyh0Fwx9B5a/
bWfUc84vv8RExnqaSF0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L7OOXKjR2mh+0VcJdUCwJQRlc+ZtxJTbvDLM2YCKpqjr0+LPmsMtcLDyB/gc14Ado9LBSJ0oay9X
3mqOuHh3uz0RTqbMOVKzN46zftuKBuzthzLrJewlP1PTtG5xH2e/VJ2QCFzTc9XsxOjW7vUt9JRf
JNwmNaVHzBkxzAEP/+z+oT2IqITTR5HWFJGKmvOFBAH8i4rPYWDmgSKN/EitHkMpEt0kSMDp3HF7
6QOkNO2ArG4aKp2yH9UEL5xHWF+fOvb1Xx9ua3KsUtuI7WeMiicZaG8uULiF5CPrytryTxYUgKbc
j/VDeDniGcP1gaQt2k86myPVyVJJz+6cPtiWPA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20672)
`protect data_block
8AOvQ/eDzj1Fhcs77c5xVvovhythjwo+rXoK4iIYXT4us9jma/pZwVEOoLDpqelaw3SUl0Cdu1Hs
adiddhFeUJ3sWPKqV03vzf2HU32iBIcSMJn2g3XZ6QM54tiZbGMwuwuShsh0ZAS1sUlolKIhUKuZ
91u06MjjwUFb03lFObU5Ym59RvWokBwJXwQCQQp9M7708XTXpVwSpGJ5jAKZATHq8sBBNaW5lhjT
3+Ylw201SBqAzkkIiEwesXEH6qQ5YphhmO/sazmVVV4kFPeEEGaVc1KJv7LpFwGdudER2rSRPw0o
uXEYIKSz1M3dp/sSDziIj2SL6kSl1eLr+gCou85Pw5BTAqpWF2dA4xgsOuSPTeBf7ud+Y1LGCOca
xTtCnzEo/g73JW4K2xY31bjV1r1Gvn4xS9B4RSVyjluNXOOl/RiF64j/7vaMDzBdEwIymVB4JAZv
WJq05O84ycwBMUKfHBptQCcTJQ4SNI2udPv/JmF9sKPnhS99zIeShxI46CIz+cKGa8g41bZsvAjN
bS7ed2Z1QVs7cM/gUJwpAyyspSr+B65WP3rXgXsAo6OJlksbK93phIH/RtB4UsOHdSpraOhP2OPD
tcqkKOO36EOBfhcVQU7BNLA96DHXtrpXUi96tVBxD8ZzGYcSau/GrhCD38sV0F/Mr3dViiOY77xJ
5HnunSuFVDixhrp3V8QOVvr1FBlcedAefyM5opBpSYOJRpb1svqoIpQ2RA0YYfWXVP6cOG+pY/0P
lZE58SzyNZh/LvbTvXKeBO8BeJWsLSFgcWVNzsWHrsJLuTYYq9mV2lF9xVOnCpnAg7gtv3KZ43kT
SwL1DSWLGtI2BzmokYOEcMBXB76s6p05/V2l5yNGclkxYjce7NdBP8XX+Nsozv85W5nUs8ER0YTZ
sSF20PsG4BqJNcGwhjeeimeE7nFp/IToLBHM83UppFA5oH4npCBFhAFwVOfwmNLkxUA2R28gCDst
F/GgVht+1hb8i5e9nRI4vBNpsp2MVRPXE0kGOk/YU7Tur9rCQMLYKx+V2rwNHQ+0r3/2y/J0er16
c1xVADxeypXRvpyK0QRkVx2qMDeFjy85qeDonWD0anHqDBiOJbn4yLK54ew/yQiHQ8ueSUcDlVfU
/FGGl8QQTAxS/e9Fcpkd6whuM791sFnIxrPEcTlqrELWY/+2K/xuTlQueSTA3mGd9MrUUvSAoAqq
ZLGnVcBhm3jxfqt2A9iX7Ak9/hrp1pMOnbjv3zXauWemsfBHkv3cnKCc9fFIso90W1PsdnuTPqDP
22O1IJ2qFrE+8UHzjKw8VMjrd8oSchC73ZsFELkMtwi3VK7MFUmI/LqYOhLJ02/bDgnLFpYcGuel
D808Pp+PHQNiA9+DPTryj1gnDSKIxwYOEO5bEHryVEAGo0jpghymIRP4pvmmoEFpZYMYfalPeTgQ
ijncmkKY9su6xmxFN4CMwA86wG2HzsB4TYCCx0WcZ6u2k1RrTsgu27To6YLvPOPMroaCsWLOJlq2
4zHU1Si/Xam1b41FAs4ekMC1APY/9U5cARA9QPPidbBnaAiIY6sYcyL3WpGSxX/IIjF1zVDsVnzG
OZHgn/bqx1CE0CKW716QDGOdU4so40lfOnxLuE4Qg0uJ1JdLXhGZ2lNtakNmcF/2uEVZoEMIsM27
kkbQ+gZVtu6av8kFY8dCaeApjHQ7KjnpvpDslyo8OIaXI1rFX48Xmv2cmCrM4es2EGpzuSMQNiw5
eSwf3P7MZlcU0vAb9oWJkkDkhzogzUjhv4BjrlXAScKcYbA3kipCZ4Hr1Vu3lRhcQfS7lIXn4KJ9
v6CrpTNwMKXo/eVcblb6UVRJC1Ie5kwurOutUneGBACS51TvzkdfVWgVTtw/FvVnWcWkqGPyKfgE
yzNUeFi9ewcbu26hVcSJeaC+gcDeNZlvnNlZ0dk7tVtsJjXRaeTs7iCLZXu7kvInfSU7Z8uIisqb
oZG5fNXa3ZXuasibeVpU+CZgyB0ibbaZf0nuS16pg5PCAD6qL1DwYTGQDOuNwhF2CsIsYdoIC6s/
gAg8p5fxdvGeXhZa8yCfvWk/CxJTVWy37lHe64OB1Hi5FxYgqSFpPz8xJcIvELQUFvzbsjbr4Kz1
szykFnV2KPTmbqIrHbWhhqSVb9KbbHYk/tyXzvoX3JoXMXRfeXWNlXqf/H6WCQTgVgTT6SIUeXcT
Wa0a6YzJIUVAYJ9kKx1b5i0CEV8gs71isozfq5Hq4laAuej85d+gwW9v2HJZ2g8X92d04MtGMwzH
6S4dcqNoIBmKRuvb4XF3gd2IFislOwVDavDjswuIvasYkaSyfLs64Uc+c6/y6meMtkmQJ5qku5Hk
aqwe5gQdULCaHuz4kEsFuHY6NihX/UyjQdYr0E0E2m8XAP0FJR9as0naTac/jrw8AqoAVPJHy8si
WaSho3OOSR9f8R/Fseg7GeGqtjHpvj14z20lpkIGQhI6m7emO0PDLz6jnlP6IfyAgKfhhYYnCqNE
soM8/EUO9XU5J1asUJi/E4q5KfCGlMvjAPzo3sGp7Ab8wtJgM08fHjfoJ6xS1fykzlzLqDAX03DF
KD2PNz32+7zMAqNeoQ9l4DJZr991Ew7Zlm27Psg6v/yrPnoBoLVydaAUQMetq+dgk7rRLDAv8K7i
OegYQellvcNL2pgO4myXatBbj94QO5p+Kxo6UaBXLDwfVKQTC9zwXWskG5LLb1IDd8aAWMThLwng
xKT1rfo6+OUkSm23udHSX5rECPcvdNSsFLEsH6Ypbz/Nhg4XjGgNYM8GW5Vrv+rzDvKTrdj1MRw8
smedXWNdg3O/FJ8ob+gagcC+YchHDbawSf67NwEsVhNWO+qZ8Ud3Czhv0IdXzOnn2wz/TxAa2BMd
h33YghiuvmPhthldA3lR+vpfgnPW56vMaGSSS9OAVqhChIRNWKSRJ5ph/z/jrtqLUqsRj8a16q6p
Cpz6BpONBzUPdNm3AK4DSMUBlofAAO4OiZWkovFOoFjDEzfMlg70g9Km263nGLuq3Phq+e6f6gpd
cBQN75r6eOEytXKjm9rEomZmZK8yscVBwdkFKhBFW5A+QIbSnV71YLt68aDgv/fCq6zbjZ6gToSx
act2+Thwn1SJPqcfp0CVzxid6KntW2CXdnn2Uoxq84MVSI9DAkFtnlKHa3J9UhBy39NOSm70lVA+
2mpBdvSka5q9MbHaAWpT65erdhnGwjZ65q6yPDOsOoMjj3u5ySgaowZwHBo/kZedsby0k8fI94dz
jQEdxoDPYb/GD1tYbL220nv5arJqN47/V/n4WUnPs90O4q/lox2THXAspb/nDNweUtRb7n3MEYQw
DPUn9fM/+vJbUw7w5n/pd8YphWX4Vl+sdP0oBuOLh3k2uooB2ctliafdZQ1lhTde5vlKi9XLCK1K
VBpTX1CA6dGkTQocFHlw1Otp+Lh/AU+caJUwmOS1ckCylDMcI538nXK7ADpG070rZS7NSTih3clC
0+/boni2pFMAhtXle7RxitfgehS0kNor6ERsIEgPw6AQc7lrKEeMOmnWggC3EVKRAmyS29YN+Aer
3TEi3YC+D7MX5HGvpupbDcZvPEm216bXo7dLFTcs+pubxIt+9rneBD8k1FyUBNFy8Oc1QhOahY6N
zMqgoTWc5NSw7+vxEdcBE6XmCppxy3FkI5mNV69HOs4DzhL8RDNVgVcHfFRPZ+1PFuSz5FCsv6/B
wW+ZfmaanVxpWo5EkXdlCpaQTONV7OP2D13BM9s+wgi9pn/0/J/w5Ifh4eI/div6qNafAXe077me
2t9MzqTgJa3II7CelqzU4CqCpG/yzXdvJi46JI025YJgA7hqPaHLbh6CRhDi16/zvz9Y5QnBLY+N
zdl4j8zYgPVHEn8YB69uzgsdSHKWpwW413SQQfKXQPhtjK8LXS3X1upNOgePVubE94mgWCVenxEz
pLei5A448wPwRJ6BZLkpqoeUxPJItPN7t38HpdBVPO/FuOSd/KUsS6YQXAxgTh5yLrP/l15K6lID
wj3MTGVQHmWjt5B+xnwAYk6tmA6th2elAH1t7Pe3n0BKUWMcyTE8/BiPVCRAJ08+N/wWK7Y+ITFY
TnFV4/iB+cU6igJlQW51XsZcT9gmbklMNF8gBDVUd8hPcQbhKbU29HJMV3erO0eeH2bRWFLV2du4
svhs3vsfaTlF029J53GdFeayx6Px/AT8KO1T7SPMpqsuNAAEyXOzoizQBmehJXzMOioN5cVYDb5K
/f+cQ7D4OiLEf2rTUSn+b5ry/1OnUBdHtEdGMFpvkzg6uET4XZCwNfE1KX5yVWXa0Vje4Sm3wV5a
K2OU/pEEIfIPqsAzSUFi5znRSigKCX8sVVGpXVTMIQezglz8dl4d9n072m8H0WYI/XW7RZj5qgMC
sZyyJ8I5mZ/J0V1DQol2LRFvvXyq2Kuqe2Q4j+MWVLS+g7InOVYcWUg7rdSxHkxO0v1C4SIgSjgr
jYVd20v39DuXWxK1qo13nqlk8zZoYuivR8TaaZLRgvPm9GccLQdMmkHKI7jbX9B+gGqCjtIBuSgO
Uea+9HGsMNrj8RlN+L3bWq6xV67EE/qLURAbl1Nke+BAAlx3nzSJTJY/2wMhP16LG+oG8fmRvIfw
+nzNd9UdcqDN+Hc+W7E+7tCYKJPuaCe0pS58UisPULqeSorHWImx7Xjt4m1DaPTEZ2VUUl3AiAiv
cJMHqokYxCC4I61k/ywuv//XMY+/G2cHmkFY+GSumFIXBnJEH3BBAeTJtZvD3jYF8OomWmbWMZCU
VVx/geQo5BxJXrRQ7kMhGbbGRR+0dOFcOUWDjCV0IfgUhp+vDrZUyy5SPHnDHRS54NkWD2qx58ld
PSfxFv+lVHoGo+uJ2jYeGvIzOumBkuJNrpOI2qW0q4ijDB1axEe+LKhnHtFK+kpxCs0mBl4oTpsC
lB86xRLnfoabAvEEVvHdLGOOACn8EkMt8TbmoAUq8jjCxBQKekn+QFDwqLYPPs/xN/9Ah3Vami2m
8jgExzxj1cYVLTr2uJMqxFNNmt6KJGLZRfSTZalmT4ig6LDbeUwuYH01u9oNITCDgBYBzmxAt/bN
iLapiIsiJAsybRk8bEY4NnkOEXA6ydBj76rFScdR6uQSC749O/tvDD7SUQqGvAH9es6B+rAbRX2h
QiKw9ntOxp91BFMsHd+gt+T/8EdGmyXR+Qu7z//0wXGo4XP+9iFluq9u5H0yIBkUk1Ex51za3l8s
rfhkYcTUOLV9fadIpNx3BVgiXhNI4mjKoCai/cJ+FQrk38ac2Ftdb0Z1AdfQdB7yY870+2SXM2vH
6Y2wUrFlELa7BVCvWf49wHhQBEeFkrDNwCNA02Tt6CRkC7Iroova/8ExgZj9HhfHbEznEgo941RS
qxFDzQieDeS8Vgn0Zwr0QRbAQLmwwBijIZ3RHbOIOCe4KYWHuVuqG4mxleUVmNgzzlgjavBpQH2M
KsgjtTElsPVFS8WSzSjSJQWBHmQJ07FFMw3tLXvtmXBMkotM8a1iqePdcFwmgz3EYv/clqct7ZwY
w9D9bocQPbHku66po3I/JD/92tbTc9tI2xaUzQR3XsyRgaIgkFFYvoYfUyGeb/cNYwYEklGoSEV4
SIGCFC2m/5MsYYp5aYzgNbKHBggtPveDHM89dAbDv6oS0IUYSYu4CqvOerJx50ShPCsanlnJq2vI
SwBREbDzw2ah+CAYe06O7YCoaUkfgcte9uDLs+aWvKnYbx3Q6daJAcgcUvI1N1djnwb6v1ZUWtbV
qeHWZtzNfORYYuFwZge2MxwY5OKL8TRXpcjjvThG64HkK7VKTRdukPo1dyp0Ub2SkCN0NQf6bkR/
zd94LARdlaJxP6I8OyjW6iGjAmg2ZBQGpDHgCx5Fek+/nAVYpx8EdXSOHrcdz4UE2lsQfT9PXB47
lnDliv2V6vfDeXIiuZ0p6Xp63C4H5aUfUMm0fClVkIubwNmZmi/bodnNrQB1ANcTiutmrdRx5zKB
lM/SU3OCYPH1E+ozLZDI7usHeFGeAF2bH1TfnxUWu3T/0XIlbZSdR+xbnxc+N7nWxfLDuRQixI7k
9QylD9ZreEsmWNiR8tRESihelKi3EAaNJiee6Byj7g6m/YKZ12Hz9N4Z5Z0ag5of7oSVhxYK0qzA
Eeh4se7eIDnUTtNLY/uxXuWKgoyj6Fv+5dhnrcbp7G2rGTc+K0R8UoF/Kmvc6GRntjvLlXFqDyfb
vO3IA5e6GAn9lGa+IFcAzmiQvUxOZ/AjKoY6v9PyHYuhB0to9X60rTm0PEqTbq7ezgu2nlYwy1TC
XWHLwdDCjCmvlcI8fteKC1L20Sky2y4IEqTEb2X7YWFNlbLiGgnlviyySa4UpercQMZOgqRbBHC4
UFyY1vTgtYc9iaoSRqzlX+gTUY1BfCGBpx2Mpr+nbYmTMzXozKVfln7drOV8aspPvRTk04vG8rsy
AtLZfsxOHAwj4y8N1u99dVngInnPFMoCRVFzK4UKUNem8pr4PQWoib8EDQ4uhq0/wCcJnp1KQLvE
E9tjBpeEPJBMs+pyJ7ALIhmBje67GuQkcxI5pEMVMvIE05gvhoH7kz4dEL+xK4Tno2z0aCitmX6K
GEzQupS1/Z/rdxuXLLzRE47ZHR68JVfXFNUsvXk0J4WZgsZDlFxRZaJbdzCgMS3xBIyIT8UCcT8S
lTZ7OGpqSfaEuR+mvAbruPG9uWPiEodtsZf3DnWkjREX0jRIMstTmLV1T/1JFtp+U3YJPS9HT+tg
/aF8NkEBpEv5gN1EK+gv7EvoKsFWtEwpfboUeOkVKPOlICG/bMW7kGkBzrCaaQg1uIOHNWLrhZQ5
NAOS8vZuzEctYOkLgx4r0yTfelt1OKH9rdcbImfOVaPYNrjHWELeeHhJ8RoHkefsD8HEmTGLkJkF
TQwC5q93SkPtMtUcJPY9uTLgAdgS/8zOeLRp6dKI/B4qndXpU9kyhVLocfzSxoW/17t/3A7009UC
4np7v9Hr+88KxOp1SbWgiVAVYQvaGw4PtbCTHWhjhSjFxO+5eqp9XcGc5h2w5kkG0XHgu/ukk3xn
jZyn6J5PKZBSIeh1hsN1ZPBKhhhtgEU6oINVNQuG5pqYwq53XwVFvqAVcVOhUcIKcWSndODw4bEa
Hyrfd1vDfx+QJiLIsswVNg8ka5PGAFfBZFZwB2zNl9Lr47ckSQf706x1MMWQ0at9oKy1Phzm0DpO
/xCdJs+yFKgO4orsxKNX3dDJ0OZeVeKXIGf21OqwlUu/dI5vIrYSglM7FCsGXC4Qe/dmzGQ4ycl2
uZIGCwjWDSwVLZrTrJU+tBXYK7YXJ/UIyvE6xLrn4SoBEvCFgfZcNEdNHR+93Tr0W7877j7VqJge
RgRLdHe975/PDYvhP94dvTYZwaO2ut/waoRJa2A/zilZbqiQJnSo2YVAFOxuNeW+S1/RoPX3ZGA/
W1eh5NQWlSwB0Pvw0+GstN93kLePYi7vEZmvkzyM8vAPiaTaIshkKA+vRX3v+TFjjPYHQ85iaeob
yoewbzvNMorL2CF20dHsJ1PUDUFHplzCwR4iuzj0aVtPnynNZzUU/+MB/sxFLhXVbegIESpegjHl
jaFQXicZJ2EES967jAvtN1FB9iE+CWtR8bGcD+01J4bS/5dKXLG8Fs0ZKdkxJE6WaIgC1jVzyDbX
BOvDuufhysCMbianfW2rLgGJYKTZ0aupcwvOC0jZznvduqXbz++KMjoxyv9SIBwHqxtCKMdkG6cU
8bxA/2gAbHSAQbAK7LnU7r8o7l4F67dpYkpnEKrr9w4AcBKqCFY1R9++6s7lEOKhq/HTSNYLS+vA
PrMsxdI36eTBe8y1kcazV1vOtm9APQsZoyJ/XcoRV3WVjfkLtpHTAOYMP9JuZJSFpkiTjBccnVYI
JIqSm8CNxe1DA4DoIx0CQs1iqp/FwGP9SCX0FC5JPcTCzqOrELGS80UNdsKpaDSWXiANQQiNskyc
5mshns2PfEfgOeujPGiRlHt+pBcsrU+ykRiqyXmODyTi1v9gKr3DSLo+32/3ZUz95GEcLLL+KwED
KpStvtkIvkilFZQB7xFiMsjBV4i1oS6Vw1W59fFprpoubg+J9CGuTc9LI9mFWy1t1Xskag7yn9vV
r7kXqBVYzjocM2IJNod3Wu3dQvqt+HxXPOsSvfam1pRbWSElrh7SN3WJLvI1aPkIQtgQLL+lRFlY
4a6azWwMNug4UKUEXEDY+welR94099waUzzGygu8iP3iy7MNFbh/MyIia0ocrKcMa2bkwq+J5Ews
hRqy/+4LtLVNRn4jPOO7wWYpwhNerSADux+EAIfv2vBVCUrANDDZkaPl6mEqEfF10GcQMd1Rtz7g
Q5MjTNTD88BDoZNXbU6IXnBRndNuMN48jTE//9O0KVNUvLxJ90kXPiQHVCo9QCdrYEdAkarY9a3f
WfnYu85CnKVM8YCwcru2p2gEleWHge2oTyv/l2Btn4eK7gSOrnMif8s0BoHiEvDM9KGmXC5tmdOz
zgvRR1fXl7vulDHz5UJ3oYAR9UnFDNjBwxLNy0+HxqwMSyFIy/fE2OC7fjlB0pkthXy9FnCZ2IVC
fwDyc4e6f2i5yCBQeiXjHtqZd57zQZVePrk3pG9ce+GDtJpRepOfeVlQiV9UHqmKIy29KvTX8bKP
W+6Cjy4xiy6lbPHQ7DON89OyLVUeiVH9ynFeELbjWB5pgZpb4sN4feCy/8Z0QLVWMnmO6y5AQQTp
4j8jhOUaLxWTJnx/34EnOEt39inT/AlMLwuSSmmtKlVuAAJW51XJl16Cgbjh1qDlSH6CgjBwy6ve
eiPYZOsbDhAgNdFp1XKtOLu2XjlDExMJbEIu/rJ1rKlX1qlaekgcpD6ATV7jV5rxtumT4OOMF7Ha
aVcH+gGX0YQQJOL5ibIsoSWxKblObefqfhZ4LJ8WKBXy1nqtmHuvPrk5/UUfKoaIgyxP7KvvlAMk
SInB89oLucvBddVImSYIdJ1svw8/hvyxKAk+JB1eqKCOKGMGxczPKTZA1+3u5mZ7a3e5MuT1d73f
ByJ/rHXTE5HNRkjdO12YS8ySPkq8Ll8MCbBwV2jMSrqPNtljBU7yydSa47uCgeCa+ozkhv/WguuY
hoK651oQwLBLL3DTfyP6urDmyVXgwHxVGGMzYC6U5husR76qb3I9xU1P1v4QBLv8i5TtDp/N6riI
r40YH18FZwVxhZUXa+huWBpsrdOZ4BwQ4BEHII8+qf7snrevQmx9Gip4iF2uYuxrMdN8GQK7wmA5
EjoIlNl9e8URGu/xzrOMWjVppaFHCz2lNuYA286FE3BYnfps56MKxVNrOeUEqqo5ptbDK48O6ETs
YqqUn4ZptprgRGs0V5nlvSdOYX2A7as8bZQF0Okdl1uoKV0PZSXmHSBTlphvgQZl5+/HXhBX53/K
lhxpV7kbKwHBBh0js8LEr3aNAzodQSMpfWD2/6GisW+gg8izWufJ4WvctTke82uup/Xv8iWdrNYu
m4tDn04zaGBTY9XxaCI4eijIryyhn7GHakHqugxpeDa5Z1MyCerrOahvEQipaCMCmMgenW89qXKy
f1K9nksDXdvrMLJOddrPpDw/EL99VhwHF8ycilgQfYyiqxZj1h8lpM8VdogIfG+m70a/yDPyMvAu
siMC4Z32I5V8WUgJvY/X9RwPZVRKH4X3HEFE22ilgsL4j3WhEC1vaYZGoy/4Z51OC4fTSIUD5/f5
IurrgDa86ekUGBpDKEx+ZBWvxfpWfO1wux1CmdxwGcnrGZ4pb+lAy+JgbaT7pjw4jQDp2GswqdTf
f1Y83lY8+qvWgb8NeWB5JMD2Qol9vd5sR+gHwhJK7abh1UBx61PfzgD4k4aMbPJkih1ia0zeuJKZ
OCtXmXlPB5Zvd0ytryJkzP2F/dRNgKlfeSHbX3k/IhswYXINLWrpi1yZxpxVyaYVyo7dAWPUGeNW
PihQQskolRWTUJTvl3jW8sr4W0ht3xLB6kxS4ICTZbNvkHOxOpZKmOP86LAJOMkA6YmYdjpyq7QM
JRczsdtxs/FrKxziY5OfX+0byJXE8id8Y82XZVat8CaF+UNKGnoFdtJGva2ts2RuHXuOC+l09ear
HyLgvAI3LJyhrWSmrgAnnR9MCDobtOPKgumm0OlbJ6/M23hBIkKMVvqoxe5I0ppI+egBsF5uwWp6
B5BzdEHspGDottMI+75W5wA4J7QNDs9NkT/2bPbGdmo1SFYe2UUWRFhnytx+mLzMzISOHyxQJ5Bm
C4FzAS4XlYp2MWzUExajQ9NHeMTz9gopbxoOLlH6PqC4Wi6UFQiQX4CJMU0FLni/Gsy8FNkxGA9y
9jZdzajdfC+8J/gccyS0xV5epVI3bPXn5zOJanPU/VuYZdSO4vLqF+Wz65v7xkcFN5eJwqvpj5i6
K0wkSlDUIdk/2NEyfppDagSgVeuii4Gi5vR+G8eMc/PGJDpuaHVP8zcT0+Tdk2P099VgEoiw9tkQ
rQ8Ecm/RB0WaHDU2r8tn8Y8TJ8LPCCq6jZozK5O8bAwTL4j0JLCoQBv9EfBxZKfbe418SIWobPiU
Vs7W8xI3afAJlEw6wzExLIch0D3INXl2Gp1mPwT+biH0xtTXgwt2GD9qmVo7gTgLSa7QvtOCxlko
Xd4ZkXA3wBnNzljgGkzjSvMTH3iAM+NTaET06xxK/zZ/5AYCQTvFCnBeJ/1bPoOB/EbjI2GVUdvT
9ntA03hb8+TP8+ZJ8TCqekp+yPRpT3KmMdQL1QWALP1UJR4Pi2IAng7CoguXpgUS5CCLyGg74Ldm
Ty+/l/l3s+T5IGLEas58p/ELwV5x+5SeyWAZILFyWemXSsmEdhOGoDbHN/A0w+MKkgPr0JBMlXBK
86aJkrvu46WFIcVErvtrg2t32JkgpWtTJa5DHrK0yL+HAvqjHrFY/BArik/kKAyRQieP4xOiHz+a
bUERwq0saacp9RX17xk131e76/RzAvujherLngbwGPagAHWeO523h10uOayBRx1aq2WQET0pOkNT
NWh6gOlk9wC4w6caWyU1Uzpq5KWwP2uMPgTCBIbtoUcOCNIbexNX5drFeGF3gRxtVpPIA71S3/v0
4xj1NdelDa2C+SjJvpgHZe5MqXKKjiFrtRTLmYY2YsZYpo97s/Z6kdkYyEO/D4TKtMStwUlu7u2k
jNiLCGmvtVUs+tg7/z7/a9WeV+Q0LddHTsE39amGJaYml4zTmKeErOzff5uuAabrq4mT4+cjJQqD
CvrYnHHzbdNvzDiv7Vx6B2xtkgPV41UBpkx5mxqoZfz8itG9D8zYlKO5uW5VTY8UTrS2lQBTrxMz
OI2COXwGVE6bARfXncPjJtag60aMb59Fl5qzXTKP9D/acbW9l40Qna5QQBP5MooaDc6NuhEsMziJ
oJbPakMlfr1p6RdMu/wNSQTgvKXiCDQ0t6wws5+sJzAHTCF876zWgUUd2iWwB/KlWUIZF1HsDmmH
LRrfn3EH2VxN+/iIRk0Gf821Hky7qdiXGPgGjp9IVbzQ66xwfXSBHfPEfACJAiU2+uqdGBX8rTxK
JKut2+zIGCjJ9GPM26A+wWDyeFiQUH50eep/FY+yINvM68+m1OVkZPPzdOYCWLyYV4OKpBLDo5hV
HXm2BtYDdlQ40VfwbWG3BB2BXxDwhvnq7aDRDbUwNlSl4CfAxP/zDueg3G00D487O+HUS+nd+o8i
o2LjfTVlShMjinyNuFIYklT+rBXGYSFU96cJbULDOA+cedT4YLi40uhVs1+QiCdNt5TVJIfjN94N
+4H5Sbb81dqZt/HaAD63WC9g5A/wIWN7npItwLfoPzhjmi/4awCtpIDBYUmV9A8PXISqQmuq99VQ
IWqzb/8vtuiJe56c3yQ4VJPg6C3pVkAy5Rk6O8+/qpScfGmx8ZwfcUQDtQ2C+8l/UEPux9FN6Big
hBGdu6UV05e1NpEds0GVDIF98ln5K5nrfeN6f9xSHuKMe2LKFp55lpUbh4CH13ak12WSLwh9Jcb7
FiFuV9w23KY6hmXrTAYXU7GE+jgX+FeA4jQbLG/ip8jUbqfkGLjNFWnfKfyP7RVMSBC3ixb5Ccz8
P+HvAN5ijPXbQfPc3GfP2cZEZ3F9rkRgF/czcqRrr1gjNZ+zFULaL5rKd8VrnadOyKlrevLQdLXq
6qzr+BTtKwcTGF7+TbJPdjGcwM3v4H/snVuqgR4JlcAFl45P34gdtxz7foKK58tSUq2N2e9wBk0c
uCE+TOV7qLHZa+aO/huanBTMsHUMjmioO/TW+WbhThBFn45M2Y/zIs0mYAzgr9s2sH2Kw3Qi5aZ2
z/nR4d4+k6jPfR3eQP2ytUPfdbJJIg6rz673d+mZG0gFb5fl2+PplrOpEZg39LIElRceT4TJSR9e
R4Ck4sYAsBbi8dhVMru/AvW8KuSbjpZpWQrQPQ/slBaGwJWx1I3eZ81cDEnurB5yzYgq340tn/CD
paTKPSrpmUS5L3pTLSJ6K2u5vmGxL6JX0J0EN1YOlKmIy5SAS9r8JecdC2NhzfZsOGtLz3EoVODJ
37VzInHnK1FJsoMN/9OQ857MOUereZZuL/UqFAJRxiLPznKyxv8wNuz35JGvt/YqyhqZRdut5tJE
wEDuomkYCzYaCZNahV37qBDNNCu2ENFf5o43dIceU5Eq+a9PsFHNVc6tv/QUDQQ2dg7IZlogA7lQ
pYXa8kuLaS96vg0/S12IRuHM3lfhZRWluqKvQeGmFuEeWv87eOONoJKSTiFcA+bOjLiLElrwie+w
ziq/ZoneqAgGm0Ye0MyMVgcSum6mQsGVWCE/YRg7KZbHzr79csiznQ5pCOrfR4WWUdqa7y/sEGdS
yj6o8gHwejcJDyhIOZO0/p9OnLWOIOfex26SeCOO1RjcyPRYwRpeuh1CMiXZ7M/kXa1ClQDzVFsY
sixpzqHTWI1KonzcheDrbfS54+dYwDdG6i663qcqTrWaLidL+qpLUZA60ENU0CLEEHgKkSkXevQw
T18PphG2M0j8Zl+QvN5nilev0QOtOQTk6hwYcasdaHnnchOHMl7SmVOXI6AhXmLqb90jLbxjlmMl
uzT7pD3Zo5vQv7MsdcBbaU3jyULANodYAZijALpVxWIUg9wmGEA9w+ZWciLoKIisK0JplqZXXJeT
xDqCXZB/Gg9R8GooVWM+Hu07SD/3xjAUmvXm6rWHFFtUgaIsGWn6UnYDyPTFGj2Q3VJejkCQV/WL
mlN1Q/mEjbLZPmNKZOdiPQCL/N9e11cpRngJIEb4k50ohg9X3pwz8ROoU/eMsluXAVWLikPE2VyN
i8Ed1m2ecEQ2KMG7pzYCEgrDuY9surokB0OgsLbvqfrLJeoHriTef+HDyISVHK430lqhyETlVS0c
kU1w5N04MK3GYbAR7aFueGiyOGJaC1kFaJZdC1UFiIFu8SaKEYKt+RdVzF6lensUOxXrcLPknKbI
83P9bmWx95tqI5yKz63J4o4yqihkyWonD4u7dT9gUZW/H9b+oZMAFEHZX+/qya4eNZLk5iY0yIp5
IKWC1lduL+UxCa4U8f1pYi44DPoFSlMg7R5yIutERnPwVPyiHzfpV/YxAx6LUAD7vqPZCxtTsVl1
SRvEPXjnL8EDF/zICJEMuAPenXSEQmxPnKTx2z8y+ZOzw+PrZ3QWv5BSo47fDvA9gsMOFSTXzhav
qG3yY2Mby9ibmXFxp6vcpRfhGGRKwcjfvUjHSJbaEnCG1CzCVBgU94UOUUvjheAISutQ2NvmyAIP
i/hR9qSIoqZVhffxsGOOL2z+yxyOWJAMS5Kh76+BJKRA/wiLW3ii2FGwz+aTmHp0a5l+sLS+1ddA
oKRGz79OvUv9KjxX0XITz4Vocqt7FvICyK0kTGPZGirysSzBEQ3wNLFoAun4AcmnB4jLssiAFfaf
NWTkGe+oAiTSd6JJ0MYQA2EI+TITg9h9SK4i6iF/uersKhuZ7NFBJupaHC8ZhcfPyj1VXCDHweK8
EKQ+y17USBL/rtgGOXA+0dcsDSn259NsoiQgP1/RSeCBJaf00BXIdCBZ+fEArymxzqHnbvICABqA
wzB01h2hMCqmLqWFccHFV2JA9+b76GIRipQB/WQuMm+M8fVFT41OuwFUV/udakJ6QBXj7PZtVWsB
lFfPJtrujvpYLZ6Fsmxh0IcIMg8nF1+ZvEmFF+6jypOb3Op9VYQSwIscyWoEUCnOo8wTGiMLkwzm
JErnhEok6ZmRYIfEhHvHx0B7gx6EEkXTYP3jhxBXxs7mfJ0uZ6UBm/UWTNB15dFWbDd255kabn3z
PMBTxTXgl0yRVBA9muGsjZdlqYD7+AaqiIx3GHXFmjt4QL+DIDlnND3V7bsu4VGdZYypufn08tlX
BxFJcDTLaJtSujRXD+7ZbQErIKLeb32SKnQVlsgocaEEtrFwLOxcI2CI6yDMK1EdvM/DJ9p5UbLn
NlWz5DR6hmjEmr3Jj7/F3ib4tfQtW+DbagRU5NSjbJT2kPijWFwY2f7GSDFALNLo9tNV8hyLpvPW
zKAQySHRdZTw/EDUA0OiqkEb0o08+XHJ/O7VV6zsPt2AgNtFNGFnnqV7kdTME6WhN1mS8pvh5cpS
cmAV0WCyLdHacdfr8WmtgM1h2OXn86uBvpT1Zbom26J9t019bC1zdr/isXVvHC5LqsAzkDQ6v4TC
1jeynp/iHbpwQbc0omaxcGaA3/Qf9lJR6YUSfK1Q15L/5Fhjhh3fVJZIT4ODy7RlJm1GyNXxdbhp
Rwbz8lAeeuiguWX35F3NSdBXKsbdVwLZUOuUoxChyXosf6a7bDIQT4lQBjDOwvcA1fGmJrRehIoU
viibpO2ObMBlzEv5Y46wuoySY3FyB3LDCzWyb8qwMzTqbE/1+8vUeFvDDH+izl2QVJD/nMdVT0U5
Q1odXRkezk5xFJQTMOubo802kB9G4kAALRRs9nhOBh/DiIDVuZWhKeUlb+pxy1yZ7cqmIG++d2zP
3KJgGBo/Y43m+1vQi94jALHx3/cjjjTFe2C+ILZnx11e93in2L/NArYwhoDBPl0w/panFHelyWs8
Bk5QXoHhAzDEuJn99iBO3znp2/wa9lyRSd5Z2kaAkcgK9PMEdlJV/zysKoF7qdZvUeMUq+yQlLrA
Ygpu8E4vjcMTAkzymgrOCMh/yNeGYodoIWuH/WFwMMOTOkkbqccYLJTzvt18lh3+/lnczO0bDdFs
GONF9C73fDxEw5l+a2u/YPFTEmC2wicw6uBWeaS/YArDNfwX9D4ep7TrIrKBONHYn0HX7bc18TJO
3LVMCjn8Sp4Up/znEGYlDzE8K4XCW9pFWnZUcLDbh0TAXLluohZEcwala9SuRQkGhmB4hlWOLfnk
J0H7kIAgNByc/044XweHIsbjsz6JzZ1r8W3G1jd6+rJwbdF5OiQJVtxFDl4R+YCqYY9hKfyLuo0c
q3nG5Q8GvwFw0LCsGW3CflowBDdcmBAB5ftEB1Cmy+wE7RJHPrJ308opXP1lLn4bmppWy2VliKi3
5gbS4BMLTRzg8ZgKMIzGziCux/Xc4Ee44zZp4LTDnazuI+i9H+68M3oJPwkld+lz48dgUpXKlhXj
N3jv8u/+b0/6elCf8SJMrEviVF47N8xALBBDEed/C9WlQcpKo2be26xgvs96+tZ20rbPTBPsl6Pa
cBvkO84Gvz0+aBFkya3zz2IdYltURGNbMxCVLi8/ZkvmUuVvb0peJA7cn+pffPbIw0moD5s1uiGR
TD2oHn2jO/avDkWqMAUEInjZpHQK1jcalZfCiPmyvPsw2SYJXuc0Kpo/nyiHenr2rhAiWZn00Mqo
dDAnmBZ8lvM9TN0Ldsdks5ATZW6yhqyMouNO5XMD6balHL8w/vPGDJoEl3MU+KKcknQ6G3U3WugC
tZ8sJ6msrQLEZmbMU2bEAlr0ayCDpAmcjKKdYIAsvxoAskSPCTyMNKiXKghCDIwdZ8IAnhRn6xA/
b4HjMuvBpUvgz8bs7rWIxiAa2/xlq1nZ8cc+PwrHO1mNpYVA2x8gyRKGm77GDpYIYbnyDSAZo2Hk
JMfBFTeIH5kqGSCA3WeIfdVc8/HQXvklNdgq5M+QK1iziYi0bqQofdrn3ot3NKVk8NEKeOzRVswJ
WWIOa/nbUP68yBw3uGDvKG/yCl62V9SkkRDO5xsfpxhMj1JtmuuCQ2X1omIqTlILNqg8RCEozpCQ
3DQij5UwJliCpa5Q8bjurg49CsgNnvtsqvOG68I5pDnoDyom0Vrh/6CWdgEoL9V3s3kKf2L2ycVv
Pbqwe6xJrLc9BMbRJlPP1jPPouRX9zp5WmyNf59oSj7Z8uaN1wRqG5ZnDpBMJuvjKX0Na86gTbJG
SQaeLXgk2epOp4RBz5QwDoIX8tnxbL0hzihDC8O1nYhQeRw7RmD3s/Ddz24mL/79jjQN2L87WpnV
7BbrhXxAsFaq1EpE9HmMOlqR0BrmVtDZmPhyBweAjNjKpbsmmRyf2riR0Yxql2xJrwjlxaJ+0Kra
6sdhU2a4HXB84FU/u08drT19rDD/9nvxHbEyzuHhDaQHk8rdRHtF2OAnEWr2X5yZuBRl6pRzKhSB
wJurfFlXDYfZoocqwsiqpNmyHwxrDLTPIhOSK58rUkZs9A9Oj01el6+ZflCcdLllKXO+kjKHADz7
t8ShHPLQnF+1vIQT+UYTt9cUuoTo4V+/Fq+xKU1Px2kkBcPmyR7SERGFgPfxmqXjZHV9j7eZHEhl
zTLWvjRHuamzRKsoCKSwDPGcdU97YKl7mH2MK74G6WtNp8h1aLNwTz5bqPWYI8RARDKSTkArAyqF
gFbhhm9Hdz7onZl/sxXpeUd8BZsEjaYiitFsgAOCMharCSdmlCMsCkxBb1Ns+5UwI+az2NzEvhR0
QQ25TBEZdrJKYWwoDjC8R9lp1tBLrRKlE+wP+IAGpNnIeP/lQ62CGlcS7EjdPARFHsV7eBru2i0d
9jYVaC2Grq/sYDdzjRGWDl3DTIRP8vhoyoGjZuEhGHN0LDkeexxXAVllYK+Gr4evO/wE1WAPmYzf
aHnjmIkOdbLNE2qpsc9FyIgMs0hE7S0tmOoJLE6xYBh1QQfpHJSOPA5bVBrkCr3kD4EuuXV37qpj
wMjOtzSMiHI1xeGjLVqT6pwAQD1U2XigFeTwoRbxS32gLmq1MIq9LN19/YbAmmLmUu6jSzpNKbsS
U5rwdPBv1g/wEtLsa6BKA2k41oN0X7+LaXSMttOsZ+Qhb71UFo4rBUdbTzBHjE3trzQn4fWZfo6Q
JAe0VLZr2iiJJ6ncYwKzgvXvIuVzmHt2Pa8H6DNXbY3ekxnz2scg+NtkWc69X9a5lgWGBLDcltd9
LDh3659VNhj6jeque7CEtGHtbYlcTtQ5lLo4ZKzbzY83uC1Ty2eaiphl/Vz54I0oOq/GkpeK5+Go
lkz7QOmbFMtPcQEHdRt1g1e7xM9mKWOHrMPpneVJdLZdS1OyoxmPX3wPu7P3m9pVsJ7LSl92DonP
kgf3/F9Kn2fpj2A66n012CG3VIhB6gpAnU7lee4pME7LwuAItlclRooPp5NmzKG8CEQHrJajONdx
I/3qQUVU7JVAQXgkZtO/uBBbU88jTWaNIi1wAcff6R3MblVu6NqFNsn35QA3Brbc0so9n8qjEAWn
diFg2r4PVFAvvCxhC6xVlpJnkAGxbRDu8Ms7xN0ELhabh0w3uWgOywBqoYjSLFxfwjVe1W0Eo0xg
fqf3MHjboKnIrhntVPyNtAsqELO6ZctmClH5Klef6y6Ap9+PuF87V3ikyCPzYdnPdzV7zonS761q
GyNKWt1REnPrx84qW2Zuc7SPQncP/6hMk0uuo2MYiXUppTzh4LzkpNOVeY3OiZPcHsmhmKBfjzzJ
iP76F1AARvylIsS9NgUAhhW/n4TJEve6lqvXsWxiPNoV12G6Z2Xxg1Xgxty9M1xeAsPcLL9SnIiK
H8ZQpF6h1CXbC+RXcOY5VZIU6g3ewQI3fp2TsEMVxZBafvMb6mityIgYq6b/PstBKWPz/CurQ726
ayt7pIDw+SdQDplBtKnovSHbVKsGPQvXMHFMRqTAGVDnNyqdBTWMaGs/fOY+lUdF2xQpk0dlRMhL
8ZnKaod6IJ6dCz4B8qKDyyr3cn1Dzy5/kmkeH4zKvDQG1hpVxqRjGl44im8OSoFNQlWY4nX9eXXA
OmD3efHuht2Qc4nTd+FRRhlVQMYc63P3zgIthIrsnTObYwqWxF44HGyx/5QBw5l9JkHfLwKmmYP/
NcRUpj7yZPOJoKktXOcmXWe67woq/GTI175tCXQIBnbvN8dVPEe7rIU8lVNIJ1DfYqu1mNKSuYP/
Abn8DqMaNJnaOTbbmcxfPFnOGOcgV9xZY5R/DiPoLbsr0IatE47JDmMX7d0QhYBXyghNZWDIArJx
+AhkwLwN0PlzRckd3wFJv/hdULXDJn7xLk0zbW22zQgPN6ZziuWq8bsKyB4NX/TcwRJF9UKB0OJi
IzILUHzzyA0MKvLIy182ptQ/DzcRFrY6+uus1/5IUaELPsRhXV+48trjLGQOlqUp8R/opzegprVb
MGHwJg/NhBZVkKkwnuMPAAk5zsKo7VLUf0azYH8Ta/e4EQc4GgvAHXs9vgHQcNsv0czhovZ9FIgz
0jd6y7NYYaHhCKV36n4UkavSedoJN2FT+Av/BH8kjIMRWRYAL58dTzb64YsswGD/1IbP8EEa+/np
+C5/+/iulxHMIodnppDuKv90RQoj/QS4CAZqqTNPKVq6MhYyNXRMISY5oErCjwnQKFiyqCciDK/Y
DgpDXZ7xBodEsqpqj07/EQWLuTezPS+gGYEFymkGi5SLwJe7/Sn2M/0Jy5/U/+b0pNmx3QtC1sk9
sO/3TJqK9xRH2JNMVgC5/HhBtUO6kKCDfzpYJWrMZkR/Op80JooSGM2y6OsLXAgAf/5bSowc3bCk
56urt2fg2ToQ3nUgzEjyLgIYilTbBOWsv956geazC6nietmQgsrV6S2FBabF7DF2Ux96z0jL1Dda
rhhKzwm50ObH3jEJztcePWqxXVMi+UHpYZYK7kDNE5B23py1Q7TltLW+wdy55yM0ffQKrRP299RW
ajgFKNYxaHFgdXOP2CW0rHKjCbm+z9N0OzkOyEddzFQwwNVHJ//xtkdfs4UMZTgHUAn/hHUutKR2
HGo18m2wJ6K7zuDf1YX/YKLZXZYrNfGfZxdFMNZv6imMLvlnn8UBxuEzMEmRcuw7aCfobIkSesFM
s7QI2oFw7NTS0p2E7MAMOTVqlj/LyCsRJBHjRG9+ukECgU6yT3rzRe+wx6rGz0vybVe33UkraCNf
Vcsm01c9jpE+B/XfCchtrKyd9aiT7kzc567MHFuMzDFV3SWr4SniqtTDnq7DPKZdygAplsBQcd1V
9JpRdIIkk4vHYpa3CiU7p7KnvrtUjGec8jJ/I9J6AkM4+LQLor/jjjor3NAuu8AjTV4CZpgrZOFH
1kpWUV8Ir61JaTvmoqR72jR8w7siX1Tv8PNO6z/JWLnrsuGpe+xSnLnvW3ObYG9uRLoZanreahAR
BSSR/MkPvyGsLc1OxNB3O0a2cprF+O7tLxeaq4Owxm82/B2drDvHF16RXSZpWsojSRi3pRE3Chan
vNbPE4LV0E/44Ez23hcDZELGX4d1TaB8f5bQJ9Vwdm0k3P5EBNC32Kz3VTrttcTxHH0yVXKZvyUZ
HK6unWN1IVoeGl1qK0o1R32069tbDT4VLQlWLlU6el2orKZbA2AacgToB9ZtVlSkaUwSQlr9L+aa
mtihSXlI4vvfHw/0RaNLu7rmLsiT9mIGXrCxIRF0pNMUWFtluKsJlNYSGEpk5zgaHmXsV5AE0Q51
p9ORQqtUGGNFyPKk1XR9mh+khbJIWtyqcldJVcJ4UALu4i0OLCdNtyRoevbYlrOR2jxVfXZSNK60
lKQdRyeHjUS69cbbWDsPf6oQFAbmmZQ5sGf2qrLUczVgTwvCV/yAF5n2MKTPHrznMW4WUx5B79vC
x9edbj3HZZPRfTwcanN4UYsBhlVTeK8VZwucpVI0V4977ZcZMwC2p3rDc6oOzB1ZDoqMF3+GJobi
65ICifDOJlue40AUotRFlg9djuf85rJ2510OKsXhHnu1/9J6NiysDoJN4s27nt51OKoXhRdbYfiW
2fiyowXZASeR4OrlUDzdPhmNXkjGSvXZUAESssaKi01GifS36/+VhSguKq1dQ9GuarUgeT8s7qDx
g4cEPFjXFDTqMi1SW7mXLShvKhdIbtUBZGTglhdukqQlHvuwHQ92oKKe3DE9EYrTr6nDMxEEY+FG
suhBr2HXZEaPvH3Jsp0ufVXATWcPuH+FJo0jT1JWmACk6BlgRNn3jV2Eh81YT9o+uaPi2g1MUs5b
LxPXJJb3RseWpehVInoFr5ynSAz2QCxDjV4rHMVM7LZQr7VmN+m3oUmukFriLaMLvSuyRn65JWFN
ItI8TOGFkkf0hfBv5J/JM/0/72GWnmc2ZQVs//tQnlygpVkJ4gR3GgaueDlEC5ansJtjIchSINtB
tA6A2pEZkYsUPLcFZWhPGbvzXlJOjPLaO58PNPoeokwBBnERCyiH24fv8uJJiOqoMR1fIeEGAZ2H
hnIrgxhZgHx/RWeqRqQc1SJam/Cz/tErvGtdj82Fh2H1PRBKqjPSqh6xNKzAXaI4IR+TSP4yQ4qG
BIFmfbvgyNkLvF3YT22peY4Ke7JsBcGjGgHrtg3p4VKukGbxws0madhF9NPHF7otnxnO0yWYP3GH
/9xOf1n9B2vGe8rMRzkKAYfvGj7p2efrc03Axe2+igzVW1oFN752hJr+bko3/1KGsIkkzlt71Ph8
R6RORDzKCd2krdP/HP5apqzPshkLRj2NYzo67JfYP1YMxZvjtxvzyETTRl7lryKxsSW/+NJJDhZC
gzuUotm2pcL3yNsM2XtiSGxc+jNYYn3H+hhe+rEmS78wxxkOlhBZnBh89MM48stdD59s5u61NjD7
HW7hYdgx5CSwQl5vugKTSGLm7CMpFFn3l+GI9TbdnObnnEMXA+jRDc4YMloWCnv/IM1hMfi3ZZMz
sJOQUA/5dy4XcMoGWtOkOviDvuviYS+9p4Bc/O1m9n99qlyu00hIJJqR12kILIVOUkadTbehMb47
6sMZuV8mmfpiFUKot5S8cjInLBnroiV/Pktn0VQCB3mMjYx3uW3PN78NYjNJ7auyBW2xI9VltBpR
SMvCU8wUgzAfNmOz+rMClkH7A9sZfgXpNMYkETDR8Wr1bcUrkIJWQAivhMmustSzaPZ2/8devYit
H6/bfRFS+Ieeeahr7tHwDa9YDCNVJK77TXA/ULAfjHAS1qHr9CRViTKTyhcJEdXrSEpSKLD/XDCu
s4b078U8h4OJL9IXYLx0ijmx9TY0eL56LmxmBoZjW+NWGb179623JQ/6qMDXqwu+019/9FzjHlGh
4EEyfoRgS9dB1MlHaBvtRy9AHVtfN3rmYVF7Z45LqFQLm5KuNw45sgD8NJrXvP1sGc/SRuPFx2qQ
LgPtAoIVNrvKC9Sw3mss1mSzTz+aYjuy8GBGkxHVuIXBwU9fey9LE70Qbq1ikl8447uqRbhMS9bO
k2/9ck+e5GiqjDAsY7Ayn3VTqAnlV6md9ompY34QyHn71unRUn91kbxr1BYSaRsy75a5lCLKJeii
0C/qoQ614yYpz0oLeZsJ+MsflzscLBOdZqfrWTKWfsEjsOGAls63W7J0H5o5p6iGq+BXesN/f5AN
wdo+tgnFLVqcUbPFGP12MgXH45e0Dp9cC6ABKdqfASV92/bsolosAC3b2/gfdJdhh695IDd3G735
5SPDA5Ahd8T9HXK7oqCsxcIecgZjTnB8qnedwd9PqCh6uZMNJQQcOpldjXJWbegEHtuVOhapzmX4
LgDqNpFMNCLIfl0JWu2JxgUzVymFEvVQuAn0WeSjd6R/HFV2oISme4k2L2yUx4VgUaof4yfprgv4
i2hGm5vVHjuKgotQhC3TiJzHYk+N2tmDrZdUk3310DXBDstFh1krrj6UgdVK/SNRezgdTRj0wpO1
Y7PxUQ3GsRMyDkCl7CuctbXxDfoyymeO2l1rTq5+0W/vJjVm6MPMYlXzqgm0VqCBGyIdekfaDrcd
dBAh08JgrQlOnsh1/ghPhtcnqVcyWJeQUvCwJFXWVJSPUq1NIgyIHuJIX7WG/BT5lFvnOOctinfX
cP4uD2dxsdr+D3h8J9oxZXz8gqi1jf1AqX7pMR9STDk9RVVhhKF5Kj1nZyrgfnMrMMi11MjBjcVw
TAHonGZm5U0xY6e5fTdQV51v1D7nOxMB7um0G86Nwuub8qgtCfN90quXohu73qVJSzN1BX+7BlMH
/2MIkGxzLO/vQr9bl7by3abH1NCD/RJheAA67U/H2Y8DKfOCevawkGjcqX4DYH5wt9MMfgg7ZuYI
YYkLZO3ICj1MT3/0vnkAgckLXN+XF2QcVByb00I3UEzzxMQiS90HTKD8+j99PwpqWYW4bLxWAPiY
PLookaKLD0N4MburWrfSk93ahTAXKdq7AtB1Z/ktZaZO9rperBLsaBupwcHMwhUawa6ey4lOYF0U
Co8k4MnE1txK3Et5I8h/8F1TAl1CL/hMI8W9A7nPz9VxUbjpTybhFHudxy58sibbex7cxwjoeXov
ncCOSgT765Sqlf+UyC/ZeOO6Zo64fjMU/xuiWDKLVBWRc8QxFSwkmFKxziPptV4QrtIfoahNPkoR
47C94ikPjGz4TUQMQVZIHMdM0DjFljy/lenpM0hVdX1VtkUCumZ9wj4y4ev/TOJCeH0ODVNQN+6y
OCzWruh8Z8RH91b5UabsyIEnkFCddLZ4qyBcMMdzT4xpqLFDWNDxXnOPb/UeOqLAK1uBeHniVmOt
GNHh+prgpv23EgN9UnTG5cnJXiL/AfJi1kr7ShnrXLnD9Re+drwzcas/IHXwl3H9e9UibbZMFYKe
tOeDugDvD/lEM/tVN4fJgPH8B8XknWMA8AswpsYQ14SQByFpZk7tq8cbl0e3u2fVihtVGGlu5aiB
dYnJ14E6021FCZxAXQdu9+UcQGmP9u4h3LqyJGjTtKX8udGOoMfXk/5RxukrDCbBW3orRd+4YF5K
58yQ7m1bB5uLdqWgYhrNKG6CSw++MMC2f+vk1rHVTI5kV1d0MslHf8Eh5d1+lJl8kyYSY7E3l9Cs
KNHLaHRvryWrUlnFxkp0id58OyukvY++3cleZZCqUKn7OBkYpgQp91bzX0O/XFAS0z8EXZGLuZOr
PapUmR3nu8AaAOJGI6B4l61UshKTtkZBQarSdWj2TIuwnChoVk1sJykKqcl7Tkd79aDrRWieBa3i
junlqDKtoAi8nEItCO8fch2znXl1Et6s2yTVX/js8Mzch0T8QLFjSMSZV0488vv7lCr7Jm0t1dkO
ejyHdOFgdmXTf20KHeacn4uuqMMTq5X6n+gkt3WPl63UN7zzMk8Sw+ckiWo6ooEuhT6K1Q2T4HgK
qUSyqTrOXJ5WnAGLzHddiscKHpHXqeRxdu2yoocb5nptnC2T4KvuK6C/8IVBT7RCerpmBTHg4+aO
wHUHh8u7jyVVzCzHM4wzxhFxnlKfgLE7N67HZtqFQ3ftHkLWY3zBOFVCC7gKKz6E20cR7np+eBpu
jtdMLwfSlF+9M6AKhwaZ3Sq1dhyr5kfo8yMKqMBK1CTmZDHom59Yt7X94GpbrRsfLZsw0Zyx7COi
YmjLqXFesxsmmNvANsy6unLkVg5ZJy0p9+OiNszQnK0B2r56r8oH87w/NbpXwZY7wQ+SFVGF9/O6
r8J2vBF5WNI2hWd3QBWjp0X9Ir1Mzcipv2cJIUYYUJLMNbDnFaER3GO+BXEK1TcEpWVv6Dvo4QBe
nYylqKjLPvTPhZJKSyD0JzIauAOklbxemspw+W8l5rYwDsi4qgFfFy5122d/ch+cuqeQVrD4yA1X
QpdJTllD4YL6KFvCx+9OO3LYvh/Mk7Qvqx5r7WkC8BES8f//KlfoBmLMH5Ph2c2IzHvNRCI/d5pz
RRtBSe6c9H7Cf+iFITR9MHiBOxVV0p8TY3kjDkqzfnt9Df0DHpo1esJZD/7jePkVFKr6pa7G/txQ
DixmssM5ZDaJEAWKUjmGA2dAPFTdtqrssH7ea6SZ3Bi7rEUqVUTRrnjWzufRIYr1+KEOzlj5QzQR
TmV1BvgZ8VktXGaflaqHp5KFP+njltMy9nNGASJphPeIkgigyCkbkeBp/DleB6UyHs/Fq98ZbIor
yd9CICSgvsLGe2M/qWVuIDsRy3hWtlVP783S/Qqh5iCEgdzfw8+7aaFqL+gQMbf7QkZCBlymrCPh
nqMXbJM+ATHkDREMPS0sEqOIr6tf0xf0QvLsxnYDqssiZbGeSh2hjv/wYkbW3YIzAPclO0OhLJEU
53rA7r+TrxmyZbrkn8zx77GoJFnhYDhwaJldd0S7UcqfmzGOIVxhb1L4MBjHSLSVpkLo2ds3gmrE
VCFnuw6MVDhQZ/HZq9XeUbEfvEsbEFDO8VnSYlTeYwp3fNz/hgJRu1NXOcbH913T1t7iKPl2/wah
f4s/W4j9mdzEcfPuDv2bWJcoZ0v+amys0W/8uVbRZyMJNtlklTP78dfmUZQrKbJGnIJO686hseAB
MuF6qb2w72jq8IlnngW23/oo71QdmjMDDH84EDSFWf5InMDL7QFzO1ZFgWO02BeDe+Yq+DThVFBp
NFGOnNy9q72mT9HiOrnMDOSScIIm3+BjGiFjGlwZcLm18x9hmkn5Ld4NHDc8WPAqYR6aatRYiGWV
VO5JfAQAZblpXSKu0htlBmsUzn2pdEjI5+0JyrHnFTeDesTnlF896Wr5VG/BLvd/TI7iaQBo1rTx
gYMcS37wtTgaj1XqLmoLmYaSgG4WSWTKm3XFaFOZpybSK9eeiLIn6E+1pfqKXEtL342k7cyrZvA+
XNBoZa6kDB3UHrivl9KTSECLq08uGgIShpnJw0ZL05clgTnKcChTrwjHGnaQecxfhNmw3pv6R7di
JcK1bBCTHVBHFpM+xpzhzDZtP5TTNq1wysOu2SY3mqjJ1zUJ1QaK5OwQ8JyM3fNdi0LAMSBkxai1
gPQGbQcONJANVwjfI7wgeDeH9qgPUFCpp7cHjLwkLwVPpCGs9wIJCWoK9zpnvXGjO7YO/vEK4Z8T
JmztuGeQBrcpocd+WO4DZjhltXWMGynrr9BrgyVy46JPujwaPpk7dbfXM3GOuErgD/qUPLrAgK7T
T19alD4zF3hqTE4Zo84hgOPcYyygAsU8YXoSw9bLvJZMnFdlJBrGOJvETXd5lRW75c4knQ5MPIVf
m/zkZoFyi/QgAlzNp04dFOi+tv3bAKzCwFBpTIuzAGbBk+IJ5DpQZx+R5Ud1ZCUi6i3UXKhQZHLi
ucXxQGYHMo/YbLj81XjYhJKJv/dUdicZhVzPxsObtQoztSXs6ulelx+V5rLceJJpeHDJbl7XKGIS
eQoElJvFuVm+SaGFzyCLNhXQRlP2Q7UthSfRnz2Zm+sn5JJHlBwVwkpyTdkaniURslZVqiwYjWdt
ZAQn+9yEsQ8VA7ymJb14vWVRvSmMZbjicEgSvyBtYlYAVewZUoyvA8z+5Kj8bP/h7UsNXOtHY/xp
JlMpvTrUCrftLV8RY75+0PiB255Ew5QAOwh+wPNR6tXUZb79Etyy4pIoBhfGKSJu914cStpKO69U
zKJBm5c0KkBl/y3v/pPIVccU7AWdpA5yHL+rR0k0vm9AhAZAJ+W/RmDubBKRT78cJQr+TD4U67DV
mNIwFn6kw2SZCJmBFvgvmnnxPbJWqjSaIUny8NRz4vIPzMmQZfiiQI7O8L+ncEqvgvlzrwzgOjFo
mNxRq+3Nv3nXePV1I9nSTMpaepiuuJmpZ8In9B5c8rvHz5D/1BLmQlkmMx+vxQy0SZaMEVRYsqBv
y8aB3g+UjM6SppVLHpCL3DuNTbWdn74ufG/BxOhSLb8KOFdYdatZ3zJmSasTtxN863QCs7NXW7Qe
lslGbEvGHkExUeWwHEVG4bf0c2wFJ0VSIDb7SKb+FLPhUWQ773egqj58kncR0OYXzKT1KlY44t8D
XZi8siaIujhzRwyZR5+Y9W5yze0+kBS1xCBZ7N+0UUCfGBqAaDecq7HDVYHxe5YxvPrGQCq5SIsM
AMmOOVdkwIfdOy9o0k4+bLLEy2HuHoLSUjQl9WKijYyw5WU3V8iAux4f9AwzKqRtfPimfz1tRlPo
3sxJREzIKV4cMTJcG8Rk5ELCCqEglgAFxhCwQgsihR4btnNIo9TZd6hhBD4uaVqD68Or1TTlxrFu
OlhBrdNFXIHjFNG5JWzD2udTq3kSTE7oGNBKKaZVzkHv+15lqJAnNLHtg18bA5kcTmiIbiGpm3V8
vgoBZV9XNohn1YzuIPEClhdB6/HTuiisVpKL2etgsioGTJ6FnauSoYQZ79eXJ/r4EPf8S0yKYx35
jNWZAowsqWp99jk5FwXsTKQeZFxMhkR4BbhRaVN1BqPVdSKjHY5VnaBdMgk0/pvHzicequGBkznx
t/+Hrbn/vi5/LwfDLktO9VJx4cX1God59HH0sljcU4l2os/EVQTj95/Dp3bLos24CHcvQz7r5Zoh
pRxXpBORlNtj6BmUDg/pMVcfw2hhCYL190MHAY6aGwrci4J1FWMxbegOAsYitcMTyl3LiVZIC3EV
qPOMqxCIO06rSiMwwwbGr4ZXMqd8R0rdNAJ+H2/Di1n700dPKGMrNl7T8RnjqulOEm20UrvFqING
y6RtNHW4pXr+XolcKMHRPpUTJadhP+lTgjYcYpO5xzYJ+2pUN8YGwzJU6sDRjzLkX9caon8/zfkF
5DILsIA9gwgoLOv/dymI6I/OFTjnxnu+5N3wibwByVP7V/xhGeqA3nShw6Gn2adCPAi8SpNab2GM
XHMFqmd3lIS7wenB3dzSBUCrbYNqzob2B8kjM8wIz1Bw/bPbW4u9yhv/j5lpo+Cs+hjpLsI0KvRs
fTPzovL09bOFErVRFwPsmk0iD+5Ou7MIXiasrxAiv3zmm3krDrvA52UFlo1knW5VSKLJM19FjWji
N1uopVub4v4VMI45q56n1EOpNyKV7gQs1oXIOlEgmZzp7OOoYdKzw6phKilzAeJ+2ffl0O7VyinI
VqbOBHESO9Fgo4r7jDNo9Yj6hRWlQ4KjCUxKs/ZiIzF53d2J5NZ92Pi5V9z5RZKUDZiHQwW0R2bG
KMhHxnd7w75IthYhEIHnVqQyE8/EO6kQ5mT5OhqxZJWsnuv1DEZTH7uqRuFlzFUGWPXpyKi1TXUX
b3gBdZyqqBkwD/vTrjLf4iug58Mp6sHoy+Ewk0OATeXyk1iLX5/ljV6gV4krOUCIjMqp8ecjb59q
HaTM6+8WPnNKMR0bm2h9tOxx1bv2gCLJ0iFoCNhFSBM4PUHyGmk8mtY/77sJCILywXsDm18Ds9aV
QD/NLlfb/Eqx4mdsIUlVE6FE5OLM/VSTdtLfdH9usk0hh1/OTTSdUy8XldJYOuqj2RJ+FMXk6sK+
rm+ESqI4dkUCqBOEYrbQLGDA/MhGi1/f1OEhen3Fxu6Z9UeF6d8=
`protect end_protected
