------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gth_quad_init.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module GTH_QUAD_init
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity GTH_QUAD_init is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;          -- Set to 1 for simulation
 
    STABLE_CLOCK_PERIOD                     : integer   := 16;  
        -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT0_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_RX_MMCM_RESET_OUT                   : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt0_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt0_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt0_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt0_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt0_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt0_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt1_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt1_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt1_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt1_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt1_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt1_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt1_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt2_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt2_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt2_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt2_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt2_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt2_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt2_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt3_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt3_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt3_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt3_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt3_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt3_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt3_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);


    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    gt0_gtrefclk0_common_in                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    gt0_qplllock_out                        : out  std_logic;
    gt0_qplllockdetclk_in                   : in   std_logic;
    gt0_qpllpd_in                           : in   std_logic;
    gt0_qpllreset_in                        : in   std_logic


);

end GTH_QUAD_init;
    
architecture RTL of GTH_QUAD_init is

--**************************Component Declarations*****************************


component GTH_QUAD 
generic
(
    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer   := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string    := "FALSE" -- Set to 1 to speed up sim reset

);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    GT0_DRP_BUSY_OUT                        : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt0_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt0_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt0_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt0_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxdlyen_in                          : in   std_logic;
    gt0_rxdlysreset_in                      : in   std_logic;
    gt0_rxdlysresetdone_out                 : out  std_logic;
    gt0_rxphalign_in                        : in   std_logic;
    gt0_rxphaligndone_out                   : out  std_logic;
    gt0_rxphalignen_in                      : in   std_logic;
    gt0_rxphdlyreset_in                     : in   std_logic;
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt0_rxsyncallin_in                      : in   std_logic;
    gt0_rxsyncdone_out                      : out  std_logic;
    gt0_rxsyncin_in                         : in   std_logic;
    gt0_rxsyncmode_in                       : in   std_logic;
    gt0_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt0_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt0_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt0_txdlyen_in                          : in   std_logic;
    gt0_txdlysreset_in                      : in   std_logic;
    gt0_txdlysresetdone_out                 : out  std_logic;
    gt0_txphalign_in                        : in   std_logic;
    gt0_txphaligndone_out                   : out  std_logic;
    gt0_txphalignen_in                      : in   std_logic;
    gt0_txphdlyreset_in                     : in   std_logic;
    gt0_txphinit_in                         : in   std_logic;
    gt0_txphinitdone_out                    : out  std_logic;
    gt0_txsyncallin_in                      : in   std_logic;
    gt0_txsyncdone_out                      : out  std_logic;
    gt0_txsyncin_in                         : in   std_logic;
    gt0_txsyncmode_in                       : in   std_logic;
    gt0_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    GT1_DRP_BUSY_OUT                        : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt1_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt1_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt1_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt1_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxdlyen_in                          : in   std_logic;
    gt1_rxdlysreset_in                      : in   std_logic;
    gt1_rxdlysresetdone_out                 : out  std_logic;
    gt1_rxphalign_in                        : in   std_logic;
    gt1_rxphaligndone_out                   : out  std_logic;
    gt1_rxphalignen_in                      : in   std_logic;
    gt1_rxphdlyreset_in                     : in   std_logic;
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt1_rxsyncallin_in                      : in   std_logic;
    gt1_rxsyncdone_out                      : out  std_logic;
    gt1_rxsyncin_in                         : in   std_logic;
    gt1_rxsyncmode_in                       : in   std_logic;
    gt1_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt1_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt1_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt1_txdlyen_in                          : in   std_logic;
    gt1_txdlysreset_in                      : in   std_logic;
    gt1_txdlysresetdone_out                 : out  std_logic;
    gt1_txphalign_in                        : in   std_logic;
    gt1_txphaligndone_out                   : out  std_logic;
    gt1_txphalignen_in                      : in   std_logic;
    gt1_txphdlyreset_in                     : in   std_logic;
    gt1_txphinit_in                         : in   std_logic;
    gt1_txphinitdone_out                    : out  std_logic;
    gt1_txsyncallin_in                      : in   std_logic;
    gt1_txsyncdone_out                      : out  std_logic;
    gt1_txsyncin_in                         : in   std_logic;
    gt1_txsyncmode_in                       : in   std_logic;
    gt1_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt1_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    GT2_DRP_BUSY_OUT                        : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt2_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt2_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt2_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt2_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxdlyen_in                          : in   std_logic;
    gt2_rxdlysreset_in                      : in   std_logic;
    gt2_rxdlysresetdone_out                 : out  std_logic;
    gt2_rxphalign_in                        : in   std_logic;
    gt2_rxphaligndone_out                   : out  std_logic;
    gt2_rxphalignen_in                      : in   std_logic;
    gt2_rxphdlyreset_in                     : in   std_logic;
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt2_rxsyncallin_in                      : in   std_logic;
    gt2_rxsyncdone_out                      : out  std_logic;
    gt2_rxsyncin_in                         : in   std_logic;
    gt2_rxsyncmode_in                       : in   std_logic;
    gt2_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt2_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt2_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt2_txdlyen_in                          : in   std_logic;
    gt2_txdlysreset_in                      : in   std_logic;
    gt2_txdlysresetdone_out                 : out  std_logic;
    gt2_txphalign_in                        : in   std_logic;
    gt2_txphaligndone_out                   : out  std_logic;
    gt2_txphalignen_in                      : in   std_logic;
    gt2_txphdlyreset_in                     : in   std_logic;
    gt2_txphinit_in                         : in   std_logic;
    gt2_txphinitdone_out                    : out  std_logic;
    gt2_txsyncallin_in                      : in   std_logic;
    gt2_txsyncdone_out                      : out  std_logic;
    gt2_txsyncin_in                         : in   std_logic;
    gt2_txsyncmode_in                       : in   std_logic;
    gt2_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt2_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    GT3_DRP_BUSY_OUT                        : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt3_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt3_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt3_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt3_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxdlyen_in                          : in   std_logic;
    gt3_rxdlysreset_in                      : in   std_logic;
    gt3_rxdlysresetdone_out                 : out  std_logic;
    gt3_rxphalign_in                        : in   std_logic;
    gt3_rxphaligndone_out                   : out  std_logic;
    gt3_rxphalignen_in                      : in   std_logic;
    gt3_rxphdlyreset_in                     : in   std_logic;
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt3_rxsyncallin_in                      : in   std_logic;
    gt3_rxsyncdone_out                      : out  std_logic;
    gt3_rxsyncin_in                         : in   std_logic;
    gt3_rxsyncmode_in                       : in   std_logic;
    gt3_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt3_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt3_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt3_txdlyen_in                          : in   std_logic;
    gt3_txdlysreset_in                      : in   std_logic;
    gt3_txdlysresetdone_out                 : out  std_logic;
    gt3_txphalign_in                        : in   std_logic;
    gt3_txphaligndone_out                   : out  std_logic;
    gt3_txphalignen_in                      : in   std_logic;
    gt3_txphdlyreset_in                     : in   std_logic;
    gt3_txphinit_in                         : in   std_logic;
    gt3_txphinitdone_out                    : out  std_logic;
    gt3_txsyncallin_in                      : in   std_logic;
    gt3_txsyncdone_out                      : out  std_logic;
    gt3_txsyncin_in                         : in   std_logic;
    gt3_txsyncmode_in                       : in   std_logic;
    gt3_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt3_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   

    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    gt0_gtrefclk0_common_in                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    gt0_qplllock_out                        : out  std_logic;
    gt0_qplllockdetclk_in                   : in   std_logic;
    gt0_qpllpd_in                           : in   std_logic;
    gt0_qpllrefclklost_out                  : out  std_logic;
    gt0_qpllreset_in                        : in   std_logic


);
end component;

component GTH_QUAD_TX_STARTUP_FSM
  Generic(
           GT_TYPE                  : string := "GTX";
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient              
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           TXUSERCLK                : in  STD_LOGIC;              --TXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;              --User Reset, can be pulled any time
           QPLLREFCLKLOST           : in  STD_LOGIC;              --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;              --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the CPLL of the GT
           TXRESETDONE              : in  STD_LOGIC;      
           MMCM_LOCK                : in  STD_LOGIC;      
           GTTXRESET                : out STD_LOGIC:='0';      
           MMCM_RESET               : out STD_LOGIC:='0';      
           QPLL_RESET               : out STD_LOGIC:='0';        --Reset QPLL
           CPLL_RESET               : out STD_LOGIC:='0';        --Reset CPLL
           TX_FSM_RESET_DONE        : out STD_LOGIC:='0';        --Reset-sequence has sucessfully been finished.
           TXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC:='0';
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';
           PHALIGNMENT_DONE         : in  STD_LOGIC;
           
           RETRY_COUNTER            : out  STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;

component GTH_QUAD_RX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           EQ_MODE                  : string := "DFE";
           GT_TYPE                  : string := "GTX";
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient                         
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;        --Stable Clock, either a stable clock from the PCB
                                                            --or reference-clock present at startup.
           RXUSERCLK                : in  STD_LOGIC;        --RXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;        --User Reset, can be pulled any time
           QPLLREFCLKLOST           : in  STD_LOGIC;        --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;        --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the CPLL of the GT
           RXRESETDONE              : in  STD_LOGIC;
           MMCM_LOCK                : in  STD_LOGIC;
           RECCLK_STABLE            : in  STD_LOGIC;
           RECCLK_MONITOR_RESTART   : in  STD_LOGIC;
           DATA_VALID               : in  STD_LOGIC;
           TXUSERRDY                : in  STD_LOGIC;       --TXUSERRDY from GT 
           DONT_RESET_ON_DATA_ERROR : in  STD_LOGIC;
           GTRXRESET                : out STD_LOGIC:='0';
           MMCM_RESET               : out STD_LOGIC:='0';
           QPLL_RESET               : out STD_LOGIC:='0';  --Reset QPLL (only if RX uses QPLL)
           CPLL_RESET               : out STD_LOGIC:='0';  --Reset CPLL (only if RX uses CPLL)
           RX_FSM_RESET_DONE        : out STD_LOGIC:='0';  --Reset-sequence has sucessfully been finished.
           RXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC;
           PHALIGNMENT_DONE         : in  STD_LOGIC; 
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';           
           RXDFEAGCHOLD             : out STD_LOGIC;
           RXDFELFHOLD              : out STD_LOGIC;
           RXLPMLFHOLD              : out STD_LOGIC;
           RXLPMHFHOLD              : out STD_LOGIC;
           RETRY_COUNTER            : out STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;




component GTH_QUAD_AUTO_PHASE_ALIGN     
  Generic(
           GT_TYPE                  : string := "GTX"
         );
    port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           RUN_PHALIGNMENT          : in  STD_LOGIC;              --Signal from the main Reset-FSM to run the auto phase-alignment procedure
           PHASE_ALIGNMENT_DONE     : out STD_LOGIC;              -- Auto phase-alignment performed sucessfully
           PHALIGNDONE              : in  STD_LOGIC;              --\ Phase-alignment signals from and to the
           DLYSRESET                : out STD_LOGIC;              -- |transceiver.
           DLYSRESETDONE            : in  STD_LOGIC;              --/
           RECCLKSTABLE             : in  STD_LOGIC               --/on the RX-side.
           
           );
end component;


component GTH_QUAD_TX_MANUAL_PHASE_ALIGN 
  Generic( NUMBER_OF_LANES          : integer range 1 to 32:= 4;  -- Number of lanes that are controlled using this FSM.
           MASTER_LANE_ID           : integer range 0 to 31:= 0   -- Number of the lane which is considered the master in manual phase-alignment
         );     

    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           RESET_PHALIGNMENT        : in  STD_LOGIC;
           RUN_PHALIGNMENT          : in  STD_LOGIC;
           PHASE_ALIGNMENT_DONE     : out STD_LOGIC := '0';       -- Manual phase-alignment performed sucessfully  
           TXDLYSRESET              : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           TXDLYSRESETDONE          : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           TXPHINIT                 : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           TXPHINITDONE             : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           TXPHALIGN                : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           TXPHALIGNDONE            : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           TXDLYEN                  : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0')
           );
end component;

component GTH_QUAD_RX_MANUAL_PHASE_ALIGN 
  Generic( NUMBER_OF_LANES          : integer range 1 to 32:= 4;  -- Number of lanes that are controlled using this FSM.
           MASTER_LANE_ID           : integer range 0 to 31:= 0   -- Number of the lane which is considered the master in manual phase-alignment
         );     

    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           RESET_PHALIGNMENT        : in  STD_LOGIC;
           RUN_PHALIGNMENT          : in  STD_LOGIC;
           PHASE_ALIGNMENT_DONE     : out STD_LOGIC := '0';       -- Manual phase-alignment performed sucessfully    
           RXDLYSRESET              : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           RXDLYSRESETDONE          : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           RXPHALIGN                : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0');
           RXPHALIGNDONE            : in  STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0);
           RXDLYEN                  : out STD_LOGIC_VECTOR(NUMBER_OF_LANES-1 downto 0) := (others=> '0')
           );
end component;

  function get_cdrlock_time(is_sim : in integer) return integer is
    variable lock_time: integer;
  begin
    if (is_sim = 1) then
      lock_time := 1000;
    else
      lock_time := 50000 / integer(6.4); --Typical CDR lock time is 50,000UI as per DS183
    end if;
    return lock_time;
  end function;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    constant RX_CDRLOCK_TIME      : integer := get_cdrlock_time(EXAMPLE_SIMULATION);       -- 200us
    constant WAIT_TIME_CDRLOCK    : integer := RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      -- 200 us time-out

    -------------------------- GT Wrapper Wires ------------------------------
    signal   gt0_txresetdone_i               : std_logic;
    signal   gt0_rxresetdone_i               : std_logic;
    signal   gt0_gttxreset_i                 : std_logic;
    signal   gt0_gttxreset_t                 : std_logic;
    signal   gt0_gtrxreset_i                 : std_logic;
    signal   gt0_gtrxreset_t                 : std_logic;
    signal   gt0_txuserrdy_i                 : std_logic;
    signal   gt0_txuserrdy_t                 : std_logic;
    signal   gt0_rxuserrdy_i                 : std_logic;
    signal   gt0_rxuserrdy_t                 : std_logic;

    signal   gt0_rxdfeagchold_i              : std_logic;
    signal   gt0_rxdfelfhold_i               : std_logic;
    signal   gt0_rxlpmlfhold_i               : std_logic;
    signal   gt0_rxlpmhfhold_i               : std_logic;


    signal   gt1_txresetdone_i               : std_logic;
    signal   gt1_rxresetdone_i               : std_logic;
    signal   gt1_gttxreset_i                 : std_logic;
    signal   gt1_gttxreset_t                 : std_logic;
    signal   gt1_gtrxreset_i                 : std_logic;
    signal   gt1_gtrxreset_t                 : std_logic;
    signal   gt1_txuserrdy_i                 : std_logic;
    signal   gt1_txuserrdy_t                 : std_logic;
    signal   gt1_rxuserrdy_i                 : std_logic;
    signal   gt1_rxuserrdy_t                 : std_logic;

    signal   gt1_rxdfeagchold_i              : std_logic;
    signal   gt1_rxdfelfhold_i               : std_logic;
    signal   gt1_rxlpmlfhold_i               : std_logic;
    signal   gt1_rxlpmhfhold_i               : std_logic;


    signal   gt2_txresetdone_i               : std_logic;
    signal   gt2_rxresetdone_i               : std_logic;
    signal   gt2_gttxreset_i                 : std_logic;
    signal   gt2_gttxreset_t                 : std_logic;
    signal   gt2_gtrxreset_i                 : std_logic;
    signal   gt2_gtrxreset_t                 : std_logic;
    signal   gt2_txuserrdy_i                 : std_logic;
    signal   gt2_txuserrdy_t                 : std_logic;
    signal   gt2_rxuserrdy_i                 : std_logic;
    signal   gt2_rxuserrdy_t                 : std_logic;

    signal   gt2_rxdfeagchold_i              : std_logic;
    signal   gt2_rxdfelfhold_i               : std_logic;
    signal   gt2_rxlpmlfhold_i               : std_logic;
    signal   gt2_rxlpmhfhold_i               : std_logic;


    signal   gt3_txresetdone_i               : std_logic;
    signal   gt3_rxresetdone_i               : std_logic;
    signal   gt3_gttxreset_i                 : std_logic;
    signal   gt3_gttxreset_t                 : std_logic;
    signal   gt3_gtrxreset_i                 : std_logic;
    signal   gt3_gtrxreset_t                 : std_logic;
    signal   gt3_txuserrdy_i                 : std_logic;
    signal   gt3_txuserrdy_t                 : std_logic;
    signal   gt3_rxuserrdy_i                 : std_logic;
    signal   gt3_rxuserrdy_t                 : std_logic;

    signal   gt3_rxdfeagchold_i              : std_logic;
    signal   gt3_rxdfelfhold_i               : std_logic;
    signal   gt3_rxlpmlfhold_i               : std_logic;
    signal   gt3_rxlpmhfhold_i               : std_logic;



    signal   gt0_qpllreset_i                 : std_logic;
    signal   gt0_qpllreset_t                 : std_logic;
    signal   gt0_qpllrefclklost_i            : std_logic;
    signal   gt0_qplllock_i                  : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_vcc_i                   : std_logic;
    signal   gt0_txphaligndone_i             : std_logic;
    signal   gt0_txdlysreset_i               : std_logic;
    signal   gt0_txdlysresetdone_i           : std_logic;
    signal   gt0_txphdlyreset_i              : std_logic;
    signal   gt0_txphalignen_i               : std_logic;
    signal   gt0_txdlyen_i                   : std_logic;
    signal   gt0_txphalign_i                 : std_logic;
    signal   gt0_txphinit_i                  : std_logic;
    signal   gt0_txphinitdone_i              : std_logic;
    signal   gt0_run_tx_phalignment_i        : std_logic;
    signal   gt0_rst_tx_phalignment_i        : std_logic;
    signal   gt0_tx_phalignment_done_i       : std_logic;
    signal   gt0_txsyncallin_i               : std_logic;
    signal   gt0_txsyncin_i                  : std_logic;
    signal   gt0_txsyncmode_i                : std_logic;
    signal   gt0_txsyncout_i                 : std_logic;
    signal   gt0_txsyncdone_i                : std_logic;

    signal   gt0_rxoutclk_i                  : std_logic;
    signal   gt0_recclk_stable_i             : std_logic;
    signal   gt0_rxphaligndone_i             : std_logic;
    signal   gt0_rxdlysreset_i               : std_logic;
    signal   gt0_rxdlysresetdone_i           : std_logic;
    signal   gt0_rxphdlyreset_i              : std_logic;
    signal   gt0_rxphalignen_i               : std_logic;
    signal   gt0_rxdlyen_i                   : std_logic;
    signal   gt0_rxphalign_i                 : std_logic;
    signal   gt0_run_rx_phalignment_i        : std_logic;
    signal   gt0_rst_rx_phalignment_i        : std_logic;
    signal   gt0_rx_phalignment_done_i       : std_logic;
    signal   gt0_rxsyncallin_i               : std_logic;
    signal   gt0_rxsyncin_i                  : std_logic;
    signal   gt0_rxsyncmode_i                : std_logic;
    signal   gt0_rxsyncout_i                 : std_logic;
    signal   gt0_rxsyncdone_i                : std_logic;
    signal   gt1_txphaligndone_i             : std_logic;
    signal   gt1_txdlysreset_i               : std_logic;
    signal   gt1_txdlysresetdone_i           : std_logic;
    signal   gt1_txphdlyreset_i              : std_logic;
    signal   gt1_txphalignen_i               : std_logic;
    signal   gt1_txdlyen_i                   : std_logic;
    signal   gt1_txphalign_i                 : std_logic;
    signal   gt1_txphinit_i                  : std_logic;
    signal   gt1_txphinitdone_i              : std_logic;
    signal   gt1_run_tx_phalignment_i        : std_logic;
    signal   gt1_rst_tx_phalignment_i        : std_logic;
    signal   gt1_tx_phalignment_done_i       : std_logic;
    signal   gt1_txsyncallin_i               : std_logic;
    signal   gt1_txsyncin_i                  : std_logic;
    signal   gt1_txsyncmode_i                : std_logic;
    signal   gt1_txsyncout_i                 : std_logic;
    signal   gt1_txsyncdone_i                : std_logic;

    signal   gt1_rxoutclk_i                  : std_logic;
    signal   gt1_recclk_stable_i             : std_logic;
    signal   gt1_rxphaligndone_i             : std_logic;
    signal   gt1_rxdlysreset_i               : std_logic;
    signal   gt1_rxdlysresetdone_i           : std_logic;
    signal   gt1_rxphdlyreset_i              : std_logic;
    signal   gt1_rxphalignen_i               : std_logic;
    signal   gt1_rxdlyen_i                   : std_logic;
    signal   gt1_rxphalign_i                 : std_logic;
    signal   gt1_run_rx_phalignment_i        : std_logic;
    signal   gt1_rst_rx_phalignment_i        : std_logic;
    signal   gt1_rx_phalignment_done_i       : std_logic;
    signal   gt1_rxsyncallin_i               : std_logic;
    signal   gt1_rxsyncin_i                  : std_logic;
    signal   gt1_rxsyncmode_i                : std_logic;
    signal   gt1_rxsyncout_i                 : std_logic;
    signal   gt1_rxsyncdone_i                : std_logic;
    signal   gt2_txphaligndone_i             : std_logic;
    signal   gt2_txdlysreset_i               : std_logic;
    signal   gt2_txdlysresetdone_i           : std_logic;
    signal   gt2_txphdlyreset_i              : std_logic;
    signal   gt2_txphalignen_i               : std_logic;
    signal   gt2_txdlyen_i                   : std_logic;
    signal   gt2_txphalign_i                 : std_logic;
    signal   gt2_txphinit_i                  : std_logic;
    signal   gt2_txphinitdone_i              : std_logic;
    signal   gt2_run_tx_phalignment_i        : std_logic;
    signal   gt2_rst_tx_phalignment_i        : std_logic;
    signal   gt2_tx_phalignment_done_i       : std_logic;
    signal   gt2_txsyncallin_i               : std_logic;
    signal   gt2_txsyncin_i                  : std_logic;
    signal   gt2_txsyncmode_i                : std_logic;
    signal   gt2_txsyncout_i                 : std_logic;
    signal   gt2_txsyncdone_i                : std_logic;

    signal   gt2_rxoutclk_i                  : std_logic;
    signal   gt2_recclk_stable_i             : std_logic;
    signal   gt2_rxphaligndone_i             : std_logic;
    signal   gt2_rxdlysreset_i               : std_logic;
    signal   gt2_rxdlysresetdone_i           : std_logic;
    signal   gt2_rxphdlyreset_i              : std_logic;
    signal   gt2_rxphalignen_i               : std_logic;
    signal   gt2_rxdlyen_i                   : std_logic;
    signal   gt2_rxphalign_i                 : std_logic;
    signal   gt2_run_rx_phalignment_i        : std_logic;
    signal   gt2_rst_rx_phalignment_i        : std_logic;
    signal   gt2_rx_phalignment_done_i       : std_logic;
    signal   gt2_rxsyncallin_i               : std_logic;
    signal   gt2_rxsyncin_i                  : std_logic;
    signal   gt2_rxsyncmode_i                : std_logic;
    signal   gt2_rxsyncout_i                 : std_logic;
    signal   gt2_rxsyncdone_i                : std_logic;
    signal   gt3_txphaligndone_i             : std_logic;
    signal   gt3_txdlysreset_i               : std_logic;
    signal   gt3_txdlysresetdone_i           : std_logic;
    signal   gt3_txphdlyreset_i              : std_logic;
    signal   gt3_txphalignen_i               : std_logic;
    signal   gt3_txdlyen_i                   : std_logic;
    signal   gt3_txphalign_i                 : std_logic;
    signal   gt3_txphinit_i                  : std_logic;
    signal   gt3_txphinitdone_i              : std_logic;
    signal   gt3_run_tx_phalignment_i        : std_logic;
    signal   gt3_rst_tx_phalignment_i        : std_logic;
    signal   gt3_tx_phalignment_done_i       : std_logic;
    signal   gt3_txsyncallin_i               : std_logic;
    signal   gt3_txsyncin_i                  : std_logic;
    signal   gt3_txsyncmode_i                : std_logic;
    signal   gt3_txsyncout_i                 : std_logic;
    signal   gt3_txsyncdone_i                : std_logic;

    signal   gt3_rxoutclk_i                  : std_logic;
    signal   gt3_recclk_stable_i             : std_logic;
    signal   gt3_rxphaligndone_i             : std_logic;
    signal   gt3_rxdlysreset_i               : std_logic;
    signal   gt3_rxdlysresetdone_i           : std_logic;
    signal   gt3_rxphdlyreset_i              : std_logic;
    signal   gt3_rxphalignen_i               : std_logic;
    signal   gt3_rxdlyen_i                   : std_logic;
    signal   gt3_rxphalign_i                 : std_logic;
    signal   gt3_run_rx_phalignment_i        : std_logic;
    signal   gt3_rst_rx_phalignment_i        : std_logic;
    signal   gt3_rx_phalignment_done_i       : std_logic;
    signal   gt3_rxsyncallin_i               : std_logic;
    signal   gt3_rxsyncin_i                  : std_logic;
    signal   gt3_rxsyncmode_i                : std_logic;
    signal   gt3_rxsyncout_i                 : std_logic;
    signal   gt3_rxsyncdone_i                : std_logic;



    --------------------------- TX Buffer Bypass Signals --------------------
    signal  mstr0_txsyncallin_i  :   std_logic;
    signal  U0_TXDLYEN           :   std_logic_vector(3 downto 0);
    signal  U0_TXDLYSRESET       :   std_logic_vector(3 downto 0);
    signal  U0_TXDLYSRESETDONE   :   std_logic_vector(3 downto 0);
    signal  U0_TXPHINIT          :   std_logic_vector(3 downto 0);
    signal  U0_TXPHINITDONE      :   std_logic_vector(3 downto 0);
    signal  U0_TXPHALIGN         :   std_logic_vector(3 downto 0);
    signal  U0_TXPHALIGNDONE     :   std_logic_vector(3 downto 0);
    signal  U0_run_tx_phalignment_i :   std_logic;
    signal  U0_rst_tx_phalignment_i :   std_logic;


    --------------------------- RX Buffer Bypass Signals --------------------
    signal   rxmstr0_rxsyncallin_i :   std_logic;
    signal   rxmstr1_rxsyncallin_i :   std_logic;
    signal   rxmstr2_rxsyncallin_i :   std_logic;
    signal   rxmstr3_rxsyncallin_i :   std_logic;


    signal   rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal      rx_cdrlocked                    : std_logic;


 


--**************************** Main Body of Code *******************************
begin
    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_vcc_i                                <= '1';

    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    GTH_QUAD_i : GTH_QUAD
    generic map
    (
        EXAMPLE_SIMULATION              =>      EXAMPLE_SIMULATION,
        WRAPPER_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP
    )
    port map
    (
        GT0_DRP_BUSY_OUT                =>      open,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X0Y0)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      gt0_drpaddr_in,
        gt0_drpclk_in                   =>      gt0_drpclk_in,
        gt0_drpdi_in                    =>      gt0_drpdi_in,
        gt0_drpdo_out                   =>      gt0_drpdo_out,
        gt0_drpen_in                    =>      gt0_drpen_in,
        gt0_drprdy_out                  =>      gt0_drprdy_out,
        gt0_drpwe_in                    =>      gt0_drpwe_in,
        ------------------------------- Loopback Ports -----------------------------
        gt0_loopback_in                 =>      gt0_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        gt0_rxpd_in                     =>      gt0_rxpd_in,
        gt0_txpd_in                     =>      gt0_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt0_rxcdrlock_out               =>      gt0_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_in,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gthrxn_in                   =>      gt0_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt0_rxdlyen_in                  =>      gt0_rxdlyen_i,
        gt0_rxdlysreset_in              =>      gt0_rxdlysreset_i,
        gt0_rxdlysresetdone_out         =>      gt0_rxdlysresetdone_i,
        gt0_rxphalign_in                =>      gt0_rxphalign_i,
        gt0_rxphaligndone_out           =>      gt0_rxphaligndone_i,
        gt0_rxphalignen_in              =>      gt0_rxphalignen_i,
        gt0_rxphdlyreset_in             =>      gt0_rxphdlyreset_i,
        gt0_rxphmonitor_out             =>      gt0_rxphmonitor_out,
        gt0_rxphslipmonitor_out         =>      gt0_rxphslipmonitor_out,
        gt0_rxsyncallin_in              =>      gt0_rxsyncallin_i,
        gt0_rxsyncdone_out              =>      gt0_rxsyncdone_i,
        gt0_rxsyncin_in                 =>      gt0_rxsyncin_i,
        gt0_rxsyncmode_in               =>      gt0_rxsyncmode_i,
        gt0_rxsyncout_out               =>      gt0_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt0_rxmcommaalignen_in          =>      gt0_rxmcommaalignen_in,
        gt0_rxpcommaalignen_in          =>      gt0_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt0_rxlpmhfhold_in              =>      gt0_rxlpmhfhold_i,
        gt0_rxlpmlfhold_in              =>      gt0_rxlpmlfhold_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt0_gthrxp_in                   =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt0_txpostcursor_in             =>      gt0_txpostcursor_in,
        gt0_txprecursor_in              =>      gt0_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_i,
        gt0_txuserrdy_in                =>      gt0_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                 =>      gt0_txusrclk_in,
        gt0_txusrclk2_in                =>      gt0_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt0_txdlyen_in                  =>      gt0_txdlyen_i,
        gt0_txdlysreset_in              =>      gt0_txdlysreset_i,
        gt0_txdlysresetdone_out         =>      gt0_txdlysresetdone_i,
        gt0_txphalign_in                =>      gt0_txphalign_i,
        gt0_txphaligndone_out           =>      gt0_txphaligndone_i,
        gt0_txphalignen_in              =>      gt0_txphalignen_i,
        gt0_txphdlyreset_in             =>      gt0_txphdlyreset_i,
        gt0_txphinit_in                 =>      gt0_txphinit_i,
        gt0_txphinitdone_out            =>      gt0_txphinitdone_i,
        gt0_txsyncallin_in              =>      gt0_txsyncallin_i,
        gt0_txsyncdone_out              =>      gt0_txsyncdone_i,
        gt0_txsyncin_in                 =>      gt0_txsyncin_i,
        gt0_txsyncmode_in               =>      gt0_txsyncmode_i,
        gt0_txsyncout_out               =>      gt0_txsyncout_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt0_txdiffctrl_in               =>      gt0_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                   =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gthtxn_out                  =>      gt0_gthtxn_out,
        gt0_gthtxp_out                  =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_out,
        gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_out,
        gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt0_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt0_txcharisk_in                =>      gt0_txcharisk_in,


        GT1_DRP_BUSY_OUT                =>      open,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X0Y1)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpaddr_in                  =>      gt1_drpaddr_in,
        gt1_drpclk_in                   =>      gt1_drpclk_in,
        gt1_drpdi_in                    =>      gt1_drpdi_in,
        gt1_drpdo_out                   =>      gt1_drpdo_out,
        gt1_drpen_in                    =>      gt1_drpen_in,
        gt1_drprdy_out                  =>      gt1_drprdy_out,
        gt1_drpwe_in                    =>      gt1_drpwe_in,
        ------------------------------- Loopback Ports -----------------------------
        gt1_loopback_in                 =>      gt1_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        gt1_rxpd_in                     =>      gt1_rxpd_in,
        gt1_txpd_in                     =>      gt1_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt1_rxuserrdy_in                =>      gt1_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      gt1_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt1_rxcdrlock_out               =>      gt1_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt1_rxusrclk_in,
        gt1_rxusrclk2_in                =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt1_rxdisperr_out               =>      gt1_rxdisperr_out,
        gt1_rxnotintable_out            =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gthrxn_in                   =>      gt1_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt1_rxdlyen_in                  =>      gt1_rxdlyen_i,
        gt1_rxdlysreset_in              =>      gt1_rxdlysreset_i,
        gt1_rxdlysresetdone_out         =>      gt1_rxdlysresetdone_i,
        gt1_rxphalign_in                =>      gt1_rxphalign_i,
        gt1_rxphaligndone_out           =>      gt1_rxphaligndone_i,
        gt1_rxphalignen_in              =>      gt1_rxphalignen_i,
        gt1_rxphdlyreset_in             =>      gt1_rxphdlyreset_i,
        gt1_rxphmonitor_out             =>      gt1_rxphmonitor_out,
        gt1_rxphslipmonitor_out         =>      gt1_rxphslipmonitor_out,
        gt1_rxsyncallin_in              =>      gt1_rxsyncallin_i,
        gt1_rxsyncdone_out              =>      gt1_rxsyncdone_i,
        gt1_rxsyncin_in                 =>      gt1_rxsyncin_i,
        gt1_rxsyncmode_in               =>      gt1_rxsyncmode_i,
        gt1_rxsyncout_out               =>      gt1_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt1_rxmcommaalignen_in          =>      gt1_rxmcommaalignen_in,
        gt1_rxpcommaalignen_in          =>      gt1_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt1_rxlpmhfhold_in              =>      gt1_rxlpmhfhold_i,
        gt1_rxlpmlfhold_in              =>      gt1_rxlpmlfhold_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt1_rxcharisk_out               =>      gt1_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt1_gthrxp_in                   =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt1_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt1_txpostcursor_in             =>      gt1_txpostcursor_in,
        gt1_txprecursor_in              =>      gt1_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_i,
        gt1_txuserrdy_in                =>      gt1_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txusrclk_in                 =>      gt1_txusrclk_in,
        gt1_txusrclk2_in                =>      gt1_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt1_txdlyen_in                  =>      gt1_txdlyen_i,
        gt1_txdlysreset_in              =>      gt1_txdlysreset_i,
        gt1_txdlysresetdone_out         =>      gt1_txdlysresetdone_i,
        gt1_txphalign_in                =>      gt1_txphalign_i,
        gt1_txphaligndone_out           =>      gt1_txphaligndone_i,
        gt1_txphalignen_in              =>      gt1_txphalignen_i,
        gt1_txphdlyreset_in             =>      gt1_txphdlyreset_i,
        gt1_txphinit_in                 =>      gt1_txphinit_i,
        gt1_txphinitdone_out            =>      gt1_txphinitdone_i,
        gt1_txsyncallin_in              =>      gt1_txsyncallin_i,
        gt1_txsyncdone_out              =>      gt1_txsyncdone_i,
        gt1_txsyncin_in                 =>      gt1_txsyncin_i,
        gt1_txsyncmode_in               =>      gt1_txsyncmode_i,
        gt1_txsyncout_out               =>      gt1_txsyncout_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt1_txdiffctrl_in               =>      gt1_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt1_txdata_in                   =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt1_gthtxn_out                  =>      gt1_gthtxn_out,
        gt1_gthtxp_out                  =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclk_out                =>      gt1_txoutclk_out,
        gt1_txoutclkfabric_out          =>      gt1_txoutclkfabric_out,
        gt1_txoutclkpcs_out             =>      gt1_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      gt1_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt1_txcharisk_in                =>      gt1_txcharisk_in,


        GT2_DRP_BUSY_OUT                =>      open,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X0Y2)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpaddr_in                  =>      gt2_drpaddr_in,
        gt2_drpclk_in                   =>      gt2_drpclk_in,
        gt2_drpdi_in                    =>      gt2_drpdi_in,
        gt2_drpdo_out                   =>      gt2_drpdo_out,
        gt2_drpen_in                    =>      gt2_drpen_in,
        gt2_drprdy_out                  =>      gt2_drprdy_out,
        gt2_drpwe_in                    =>      gt2_drpwe_in,
        ------------------------------- Loopback Ports -----------------------------
        gt2_loopback_in                 =>      gt2_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        gt2_rxpd_in                     =>      gt2_rxpd_in,
        gt2_txpd_in                     =>      gt2_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt2_rxuserrdy_in                =>      gt2_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      gt2_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt2_rxcdrlock_out               =>      gt2_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt2_rxusrclk_in,
        gt2_rxusrclk2_in                =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt2_rxdisperr_out               =>      gt2_rxdisperr_out,
        gt2_rxnotintable_out            =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gthrxn_in                   =>      gt2_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt2_rxdlyen_in                  =>      gt2_rxdlyen_i,
        gt2_rxdlysreset_in              =>      gt2_rxdlysreset_i,
        gt2_rxdlysresetdone_out         =>      gt2_rxdlysresetdone_i,
        gt2_rxphalign_in                =>      gt2_rxphalign_i,
        gt2_rxphaligndone_out           =>      gt2_rxphaligndone_i,
        gt2_rxphalignen_in              =>      gt2_rxphalignen_i,
        gt2_rxphdlyreset_in             =>      gt2_rxphdlyreset_i,
        gt2_rxphmonitor_out             =>      gt2_rxphmonitor_out,
        gt2_rxphslipmonitor_out         =>      gt2_rxphslipmonitor_out,
        gt2_rxsyncallin_in              =>      gt2_rxsyncallin_i,
        gt2_rxsyncdone_out              =>      gt2_rxsyncdone_i,
        gt2_rxsyncin_in                 =>      gt2_rxsyncin_i,
        gt2_rxsyncmode_in               =>      gt2_rxsyncmode_i,
        gt2_rxsyncout_out               =>      gt2_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt2_rxmcommaalignen_in          =>      gt2_rxmcommaalignen_in,
        gt2_rxpcommaalignen_in          =>      gt2_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt2_rxlpmhfhold_in              =>      gt2_rxlpmhfhold_i,
        gt2_rxlpmlfhold_in              =>      gt2_rxlpmlfhold_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt2_rxcharisk_out               =>      gt2_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt2_gthrxp_in                   =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt2_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt2_txpostcursor_in             =>      gt2_txpostcursor_in,
        gt2_txprecursor_in              =>      gt2_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_i,
        gt2_txuserrdy_in                =>      gt2_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txusrclk_in                 =>      gt2_txusrclk_in,
        gt2_txusrclk2_in                =>      gt2_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt2_txdlyen_in                  =>      gt2_txdlyen_i,
        gt2_txdlysreset_in              =>      gt2_txdlysreset_i,
        gt2_txdlysresetdone_out         =>      gt2_txdlysresetdone_i,
        gt2_txphalign_in                =>      gt2_txphalign_i,
        gt2_txphaligndone_out           =>      gt2_txphaligndone_i,
        gt2_txphalignen_in              =>      gt2_txphalignen_i,
        gt2_txphdlyreset_in             =>      gt2_txphdlyreset_i,
        gt2_txphinit_in                 =>      gt2_txphinit_i,
        gt2_txphinitdone_out            =>      gt2_txphinitdone_i,
        gt2_txsyncallin_in              =>      gt2_txsyncallin_i,
        gt2_txsyncdone_out              =>      gt2_txsyncdone_i,
        gt2_txsyncin_in                 =>      gt2_txsyncin_i,
        gt2_txsyncmode_in               =>      gt2_txsyncmode_i,
        gt2_txsyncout_out               =>      gt2_txsyncout_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt2_txdiffctrl_in               =>      gt2_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt2_txdata_in                   =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt2_gthtxn_out                  =>      gt2_gthtxn_out,
        gt2_gthtxp_out                  =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclk_out                =>      gt2_txoutclk_out,
        gt2_txoutclkfabric_out          =>      gt2_txoutclkfabric_out,
        gt2_txoutclkpcs_out             =>      gt2_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      gt2_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt2_txcharisk_in                =>      gt2_txcharisk_in,


        GT3_DRP_BUSY_OUT                =>      open,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X0Y3)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpaddr_in                  =>      gt3_drpaddr_in,
        gt3_drpclk_in                   =>      gt3_drpclk_in,
        gt3_drpdi_in                    =>      gt3_drpdi_in,
        gt3_drpdo_out                   =>      gt3_drpdo_out,
        gt3_drpen_in                    =>      gt3_drpen_in,
        gt3_drprdy_out                  =>      gt3_drprdy_out,
        gt3_drpwe_in                    =>      gt3_drpwe_in,
        ------------------------------- Loopback Ports -----------------------------
        gt3_loopback_in                 =>      gt3_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        gt3_rxpd_in                     =>      gt3_rxpd_in,
        gt3_txpd_in                     =>      gt3_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt3_rxuserrdy_in                =>      gt3_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      gt3_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt3_rxcdrlock_out               =>      gt3_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt3_rxusrclk_in,
        gt3_rxusrclk2_in                =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt3_rxdisperr_out               =>      gt3_rxdisperr_out,
        gt3_rxnotintable_out            =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gthrxn_in                   =>      gt3_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt3_rxdlyen_in                  =>      gt3_rxdlyen_i,
        gt3_rxdlysreset_in              =>      gt3_rxdlysreset_i,
        gt3_rxdlysresetdone_out         =>      gt3_rxdlysresetdone_i,
        gt3_rxphalign_in                =>      gt3_rxphalign_i,
        gt3_rxphaligndone_out           =>      gt3_rxphaligndone_i,
        gt3_rxphalignen_in              =>      gt3_rxphalignen_i,
        gt3_rxphdlyreset_in             =>      gt3_rxphdlyreset_i,
        gt3_rxphmonitor_out             =>      gt3_rxphmonitor_out,
        gt3_rxphslipmonitor_out         =>      gt3_rxphslipmonitor_out,
        gt3_rxsyncallin_in              =>      gt3_rxsyncallin_i,
        gt3_rxsyncdone_out              =>      gt3_rxsyncdone_i,
        gt3_rxsyncin_in                 =>      gt3_rxsyncin_i,
        gt3_rxsyncmode_in               =>      gt3_rxsyncmode_i,
        gt3_rxsyncout_out               =>      gt3_rxsyncout_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt3_rxmcommaalignen_in          =>      gt3_rxmcommaalignen_in,
        gt3_rxpcommaalignen_in          =>      gt3_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt3_rxlpmhfhold_in              =>      gt3_rxlpmhfhold_i,
        gt3_rxlpmlfhold_in              =>      gt3_rxlpmlfhold_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt3_rxcharisk_out               =>      gt3_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt3_gthrxp_in                   =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt3_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt3_txpostcursor_in             =>      gt3_txpostcursor_in,
        gt3_txprecursor_in              =>      gt3_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_i,
        gt3_txuserrdy_in                =>      gt3_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txusrclk_in                 =>      gt3_txusrclk_in,
        gt3_txusrclk2_in                =>      gt3_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        gt3_txdlyen_in                  =>      gt3_txdlyen_i,
        gt3_txdlysreset_in              =>      gt3_txdlysreset_i,
        gt3_txdlysresetdone_out         =>      gt3_txdlysresetdone_i,
        gt3_txphalign_in                =>      gt3_txphalign_i,
        gt3_txphaligndone_out           =>      gt3_txphaligndone_i,
        gt3_txphalignen_in              =>      gt3_txphalignen_i,
        gt3_txphdlyreset_in             =>      gt3_txphdlyreset_i,
        gt3_txphinit_in                 =>      gt3_txphinit_i,
        gt3_txphinitdone_out            =>      gt3_txphinitdone_i,
        gt3_txsyncallin_in              =>      gt3_txsyncallin_i,
        gt3_txsyncdone_out              =>      gt3_txsyncdone_i,
        gt3_txsyncin_in                 =>      gt3_txsyncin_i,
        gt3_txsyncmode_in               =>      gt3_txsyncmode_i,
        gt3_txsyncout_out               =>      gt3_txsyncout_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt3_txdiffctrl_in               =>      gt3_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt3_txdata_in                   =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt3_gthtxn_out                  =>      gt3_gthtxn_out,
        gt3_gthtxp_out                  =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclk_out                =>      gt3_txoutclk_out,
        gt3_txoutclkfabric_out          =>      gt3_txoutclkfabric_out,
        gt3_txoutclkpcs_out             =>      gt3_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      gt3_txresetdone_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt3_txcharisk_in                =>      gt3_txcharisk_in,




    --____________________________COMMON PORTS________________________________
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        gt0_gtrefclk0_common_in         =>      gt0_gtrefclk0_common_in,
        ------------------------- Common Block - QPLL Ports ------------------------
        gt0_qplllock_out                =>      gt0_qplllock_i,
        gt0_qplllockdetclk_in           =>      gt0_qplllockdetclk_in,
        gt0_qpllpd_in                   =>      gt0_qpllpd_in,
        gt0_qpllrefclklost_out          =>      gt0_qpllrefclklost_i,
        gt0_qpllreset_in                =>      gt0_qpllreset_i

    );




GT0_TXRESETDONE_OUT                          <= gt0_txresetdone_i;
GT0_RXRESETDONE_OUT                          <= gt0_rxresetdone_i;
GT0_RXOUTCLK_OUT                             <= gt0_rxoutclk_i;
GT1_TXRESETDONE_OUT                          <= gt1_txresetdone_i;
GT1_RXRESETDONE_OUT                          <= gt1_rxresetdone_i;
GT1_RXOUTCLK_OUT                             <= gt1_rxoutclk_i;
GT2_TXRESETDONE_OUT                          <= gt2_txresetdone_i;
GT2_RXRESETDONE_OUT                          <= gt2_rxresetdone_i;
GT2_RXOUTCLK_OUT                             <= gt2_rxoutclk_i;
GT3_TXRESETDONE_OUT                          <= gt3_txresetdone_i;
GT3_RXRESETDONE_OUT                          <= gt3_rxresetdone_i;
GT3_RXOUTCLK_OUT                             <= gt3_rxoutclk_i;
GT0_QPLLLOCK_OUT                             <= gt0_qplllock_i;

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    gt0_gttxreset_i                              <= GT0_GTTXRESET_IN or gt0_gttxreset_t;
    gt0_gtrxreset_i                              <= GT0_GTRXRESET_IN or gt0_gtrxreset_t;
    gt0_txuserrdy_i                              <= GT0_TXUSERRDY_IN or gt0_txuserrdy_t;
    gt0_rxuserrdy_i                              <= GT0_RXUSERRDY_IN or gt0_rxuserrdy_t;
    gt1_gttxreset_i                              <= GT1_GTTXRESET_IN or gt1_gttxreset_t;
    gt1_gtrxreset_i                              <= GT1_GTRXRESET_IN or gt1_gtrxreset_t;
    gt1_txuserrdy_i                              <= GT1_TXUSERRDY_IN or gt1_txuserrdy_t;
    gt1_rxuserrdy_i                              <= GT1_RXUSERRDY_IN or gt1_rxuserrdy_t;
    gt2_gttxreset_i                              <= GT2_GTTXRESET_IN or gt2_gttxreset_t;
    gt2_gtrxreset_i                              <= GT2_GTRXRESET_IN or gt2_gtrxreset_t;
    gt2_txuserrdy_i                              <= GT2_TXUSERRDY_IN or gt2_txuserrdy_t;
    gt2_rxuserrdy_i                              <= GT2_RXUSERRDY_IN or gt2_rxuserrdy_t;
    gt3_gttxreset_i                              <= GT3_GTTXRESET_IN or gt3_gttxreset_t;
    gt3_gtrxreset_i                              <= GT3_GTRXRESET_IN or gt3_gtrxreset_t;
    gt3_txuserrdy_i                              <= GT3_TXUSERRDY_IN or gt3_txuserrdy_t;
    gt3_rxuserrdy_i                              <= GT3_RXUSERRDY_IN or gt3_rxuserrdy_t;
    gt0_qpllreset_i                              <= GT0_QPLLRESET_IN or gt0_qpllreset_t;
end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate
gt0_gttxreset_i                              <= gt0_gttxreset_t;
gt0_gtrxreset_i                              <= gt0_gtrxreset_t;
gt0_txuserrdy_i                              <= gt0_txuserrdy_t;
gt0_rxuserrdy_i                              <= gt0_rxuserrdy_t;
gt1_gttxreset_i                              <= gt1_gttxreset_t;
gt1_gtrxreset_i                              <= gt1_gtrxreset_t;
gt1_txuserrdy_i                              <= gt1_txuserrdy_t;
gt1_rxuserrdy_i                              <= gt1_rxuserrdy_t;
gt2_gttxreset_i                              <= gt2_gttxreset_t;
gt2_gtrxreset_i                              <= gt2_gtrxreset_t;
gt2_txuserrdy_i                              <= gt2_txuserrdy_t;
gt2_rxuserrdy_i                              <= gt2_rxuserrdy_t;
gt3_gttxreset_i                              <= gt3_gttxreset_t;
gt3_gtrxreset_i                              <= gt3_gtrxreset_t;
gt3_txuserrdy_i                              <= gt3_txuserrdy_t;
gt3_rxuserrdy_i                              <= gt3_rxuserrdy_t;
gt0_qpllreset_i                              <= gt0_qpllreset_t;
end generate no_chipscope;


gt0_txresetfsm_i:  GTH_QUAD_TX_STARTUP_FSM 

  generic map(
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT0_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt0_txresetdone_i,
        MMCM_LOCK                       =>      GT0_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt0_gttxreset_t,
        MMCM_RESET                      =>      GT0_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      gt0_qpllreset_t,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT0_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt0_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt0_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt0_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt1_txresetfsm_i:  GTH_QUAD_TX_STARTUP_FSM 

  generic map(
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT1_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt1_txresetdone_i,
        MMCM_LOCK                       =>      GT1_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt1_gttxreset_t,
        MMCM_RESET                      =>      GT1_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT1_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt1_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt1_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt1_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt2_txresetfsm_i:  GTH_QUAD_TX_STARTUP_FSM 

  generic map(
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT2_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt2_txresetdone_i,
        MMCM_LOCK                       =>      GT2_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt2_gttxreset_t,
        MMCM_RESET                      =>      GT2_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT2_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt2_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt2_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt2_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );

gt3_txresetfsm_i:  GTH_QUAD_TX_STARTUP_FSM 

  generic map(
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => TRUE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT3_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        TXRESETDONE                     =>      gt3_txresetdone_i,
        MMCM_LOCK                       =>      GT3_TX_MMCM_LOCK_IN,
        GTTXRESET                       =>      gt3_gttxreset_t,
        MMCM_RESET                      =>      GT3_TX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        TX_FSM_RESET_DONE               =>      GT3_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt3_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt3_run_tx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt3_rst_tx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_tx_phalignment_done_i,
        RETRY_COUNTER                   =>      open
           );





gt0_rxresetfsm_i:  GTH_QUAD_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT0_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt0_rxresetdone_i,
        MMCM_LOCK                       =>      GT0_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT0_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt0_gtrxreset_t,
        MMCM_RESET                      =>      GT0_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT0_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt0_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt0_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt0_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt0_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt0_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt0_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt0_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt0_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );

gt1_rxresetfsm_i:  GTH_QUAD_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT1_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt1_rxresetdone_i,
        MMCM_LOCK                       =>      GT1_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt1_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT1_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt1_gtrxreset_t,
        MMCM_RESET                      =>      GT1_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT1_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt1_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt1_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt1_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt1_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt1_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt1_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt1_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt1_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );

gt2_rxresetfsm_i:  GTH_QUAD_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT2_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt2_rxresetdone_i,
        MMCM_LOCK                       =>      GT2_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt2_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT2_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt2_gtrxreset_t,
        MMCM_RESET                      =>      GT2_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT2_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt2_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt2_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt2_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt2_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt2_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt2_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt2_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt2_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );

gt3_rxresetfsm_i:  GTH_QUAD_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTH", --GTX or GTH or GTP
           EQ_MODE                  => "LPM",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => TRUE ,                        -- the TX and RX Reset FSMs must 
           RX_QPLL_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT3_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_i,
        CPLLREFCLKLOST                  =>      tied_to_ground_i,
        QPLLLOCK                        =>      gt0_qplllock_i,
        CPLLLOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt3_rxresetdone_i,
        MMCM_LOCK                       =>      GT3_RX_MMCM_LOCK_IN,
        RECCLK_STABLE                   =>      gt3_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT3_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt3_gtrxreset_t,
        MMCM_RESET                      =>      GT3_RX_MMCM_RESET_OUT,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT3_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt3_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      gt3_run_rx_phalignment_i,
        RESET_PHALIGNMENT               =>      gt3_rst_rx_phalignment_i,
        PHALIGNMENT_DONE                =>      gt3_rx_phalignment_done_i,
        RXDFEAGCHOLD                    =>      gt3_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt3_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt3_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt3_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



  cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt0_gtrxreset_i = '1') then
          rx_cdrlocked       <= '0';
          rx_cdrlock_counter <=  0                        after DLY;
        elsif (rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          rx_cdrlocked       <= '1';
          rx_cdrlock_counter <= rx_cdrlock_counter        after DLY;
        else
          rx_cdrlock_counter <= rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

gt0_recclk_stable_i                          <= rx_cdrlocked;
gt1_recclk_stable_i                          <= rx_cdrlocked;
gt2_recclk_stable_i                          <= rx_cdrlocked;
gt3_recclk_stable_i                          <= rx_cdrlocked;



    --------------------------- TX Buffer Bypass Logic --------------------
    -- The TX SYNC Module drives the ports needed to Bypass the TX Buffer.
    -- Include the TX SYNC module in your own design if TX Buffer is bypassed.

--Manual
   gt0_tx_manual_phase_i : GTH_QUAD_TX_MANUAL_PHASE_ALIGN
   generic map
   ( NUMBER_OF_LANES	  => 4,
     MASTER_LANE_ID       =>  0
   )
   port map
   (
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RESET_PHALIGNMENT               =>      U0_rst_tx_phalignment_i,   --TODO
        RUN_PHALIGNMENT                 =>      U0_run_tx_phalignment_i,      --TODO
        PHASE_ALIGNMENT_DONE            =>      gt0_tx_phalignment_done_i,
        TXDLYSRESET                     =>      U0_TXDLYSRESET,
        TXDLYSRESETDONE                 =>      U0_TXDLYSRESETDONE,
        TXPHINIT                        =>      U0_TXPHINIT,
        TXPHINITDONE                    =>      U0_TXPHINITDONE,
        TXPHALIGN                       =>      U0_TXPHALIGN,
        TXPHALIGNDONE                   =>      U0_TXPHALIGNDONE,
        TXDLYEN                         =>      U0_TXDLYEN
   );

gt0_txphdlyreset_i                           <= tied_to_ground_i;
gt0_txphalignen_i                            <= tied_to_vcc_i;
gt0_txdlysreset_i                            <= U0_TXDLYSRESET(0);
gt0_txphinit_i                               <= U0_TXPHINIT(0);
gt0_txphalign_i                              <= U0_TXPHALIGN(0);
gt0_txdlyen_i                                <= U0_TXDLYEN(0);
U0_TXDLYSRESETDONE(0)                        <= gt0_txdlysresetdone_i;
U0_TXPHINITDONE(0)                           <= gt0_txphinitdone_i;
U0_TXPHALIGNDONE(0)                          <= gt0_txphaligndone_i;

gt0_txsyncallin_i                            <= gt0_txphaligndone_i;
gt0_txsyncin_i                               <= gt0_txsyncout_i;
gt0_txsyncmode_i                             <= tied_to_vcc_i;

 
gt1_txdlysreset_i                            <= U0_TXDLYSRESET(1);
gt1_txphinit_i                               <= U0_TXPHINIT(1);
gt1_txphalign_i                              <= U0_TXPHALIGN(1);
gt1_txphalignen_i                            <= tied_to_vcc_i;
gt1_txphdlyreset_i                           <= tied_to_ground_i;
gt1_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(1)                        <= gt1_txdlysresetdone_i;
U0_TXPHINITDONE(1)                           <= gt1_txphinitdone_i;
U0_TXPHALIGNDONE(1)                          <= gt1_txphaligndone_i;

gt1_txsyncallin_i                            <= tied_to_ground_i;
gt1_txsyncin_i                               <= tied_to_ground_i;
gt1_txsyncmode_i                             <= tied_to_ground_i;
 
gt2_txdlysreset_i                            <= U0_TXDLYSRESET(2);
gt2_txphinit_i                               <= U0_TXPHINIT(2);
gt2_txphalign_i                              <= U0_TXPHALIGN(2);
gt2_txphalignen_i                            <= tied_to_vcc_i;
gt2_txphdlyreset_i                           <= tied_to_ground_i;
gt2_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(2)                        <= gt2_txdlysresetdone_i;
U0_TXPHINITDONE(2)                           <= gt2_txphinitdone_i;
U0_TXPHALIGNDONE(2)                          <= gt2_txphaligndone_i;

gt2_txsyncallin_i                            <= tied_to_ground_i;
gt2_txsyncin_i                               <= tied_to_ground_i;
gt2_txsyncmode_i                             <= tied_to_ground_i;
 
gt3_txdlysreset_i                            <= U0_TXDLYSRESET(3);
gt3_txphinit_i                               <= U0_TXPHINIT(3);
gt3_txphalign_i                              <= U0_TXPHALIGN(3);
gt3_txphalignen_i                            <= tied_to_vcc_i;
gt3_txphdlyreset_i                           <= tied_to_ground_i;
gt3_txdlyen_i                                <= tied_to_ground_i;
U0_TXDLYSRESETDONE(3)                        <= gt3_txdlysresetdone_i;
U0_TXPHINITDONE(3)                           <= gt3_txphinitdone_i;
U0_TXPHALIGNDONE(3)                          <= gt3_txphaligndone_i;

gt3_txsyncallin_i                            <= tied_to_ground_i;
gt3_txsyncin_i                               <= tied_to_ground_i;
gt3_txsyncmode_i                             <= tied_to_ground_i;

    U0_run_tx_phalignment_i    <=  gt0_run_tx_phalignment_i 
 
                                             and gt1_run_tx_phalignment_i
 
                                             and gt2_run_tx_phalignment_i
 
                                             and gt3_run_tx_phalignment_i
                                             ;

    U0_rst_tx_phalignment_i    <=  gt0_rst_tx_phalignment_i 
 
                                             or gt1_rst_tx_phalignment_i
 
                                             or gt2_rst_tx_phalignment_i
 
                                             or gt3_rst_tx_phalignment_i
                                             ;



   --------------------------- RX Buffer Bypass Logic --------------------
--   The RX SYNC Module drives the ports needed to Bypass the RX Buffer.
--   Include the RX SYNC module in your own design if RX Buffer is bypassed.


--Auto

gt0_rxphdlyreset_i                           <= tied_to_ground_i;
gt0_rxphalignen_i                            <= tied_to_ground_i;
gt0_rxdlyen_i                                <= tied_to_ground_i;
gt0_rxphalign_i                              <= tied_to_ground_i;
gt0_rxsyncallin_i                            <= gt0_rxphaligndone_i;
gt0_rxsyncin_i                               <= gt0_rxsyncout_i;
gt0_rxsyncmode_i                             <= tied_to_vcc_i;


gt0_rx_auto_phase_align_i : GTH_QUAD_AUTO_PHASE_ALIGN    
  generic map(
                 GT_TYPE                  => "GTH" --GTX or GTH or GTP
             )
  port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt0_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt0_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt0_rxsyncdone_i,
        DLYSRESET                       =>      gt0_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt0_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt0_recclk_stable_i
     );



--Auto

gt1_rxphdlyreset_i                           <= tied_to_ground_i;
gt1_rxphalignen_i                            <= tied_to_ground_i;
gt1_rxdlyen_i                                <= tied_to_ground_i;
gt1_rxphalign_i                              <= tied_to_ground_i;
gt1_rxsyncallin_i                            <= gt1_rxphaligndone_i;
gt1_rxsyncin_i                               <= gt1_rxsyncout_i;
gt1_rxsyncmode_i                             <= tied_to_vcc_i;


gt1_rx_auto_phase_align_i : GTH_QUAD_AUTO_PHASE_ALIGN    
  generic map(
                 GT_TYPE                  => "GTH" --GTX or GTH or GTP
             )
  port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt1_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt1_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt1_rxsyncdone_i,
        DLYSRESET                       =>      gt1_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt1_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt1_recclk_stable_i
     );



--Auto

gt2_rxphdlyreset_i                           <= tied_to_ground_i;
gt2_rxphalignen_i                            <= tied_to_ground_i;
gt2_rxdlyen_i                                <= tied_to_ground_i;
gt2_rxphalign_i                              <= tied_to_ground_i;
gt2_rxsyncallin_i                            <= gt2_rxphaligndone_i;
gt2_rxsyncin_i                               <= gt2_rxsyncout_i;
gt2_rxsyncmode_i                             <= tied_to_vcc_i;


gt2_rx_auto_phase_align_i : GTH_QUAD_AUTO_PHASE_ALIGN    
  generic map(
                 GT_TYPE                  => "GTH" --GTX or GTH or GTP
             )
  port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt2_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt2_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt2_rxsyncdone_i,
        DLYSRESET                       =>      gt2_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt2_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt2_recclk_stable_i
     );



--Auto

gt3_rxphdlyreset_i                           <= tied_to_ground_i;
gt3_rxphalignen_i                            <= tied_to_ground_i;
gt3_rxdlyen_i                                <= tied_to_ground_i;
gt3_rxphalign_i                              <= tied_to_ground_i;
gt3_rxsyncallin_i                            <= gt3_rxphaligndone_i;
gt3_rxsyncin_i                               <= gt3_rxsyncout_i;
gt3_rxsyncmode_i                             <= tied_to_vcc_i;


gt3_rx_auto_phase_align_i : GTH_QUAD_AUTO_PHASE_ALIGN    
  generic map(
                 GT_TYPE                  => "GTH" --GTX or GTH or GTP
             )
  port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RUN_PHALIGNMENT                 =>      gt3_run_rx_phalignment_i,
        PHASE_ALIGNMENT_DONE            =>      gt3_rx_phalignment_done_i,
        PHALIGNDONE                     =>      gt3_rxsyncdone_i,
        DLYSRESET                       =>      gt3_rxdlysreset_i,
        DLYSRESETDONE                   =>      gt3_rxdlysresetdone_i,
        RECCLKSTABLE                    =>      gt3_recclk_stable_i
     );



end RTL;


