-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : gtx_minipod_12x_k7.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gtx_minipod_12x_k7 (a GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity gtx_minipod_12x_k7 is
generic
(
    QPLL_FBDIV_TOP                 : integer  := 16;

    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP     : string     :=  "FALSE";        -- Set to "true" to speed up sim reset
    RX_DFE_KL_CFG2_IN               : bit_vector :=  X"301148AC";
    PMA_RSV_IN                      : bit_vector :=  x"00018480"

);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT0_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT0_CPLLLOCK_OUT                        : out  std_logic;
    GT0_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT0_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT0_DRPCLK_IN                           : in   std_logic;
    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT0_DRPEN_IN                            : in   std_logic;
    GT0_DRPRDY_OUT                          : out  std_logic;
    GT0_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT0_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT0_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT0_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT0_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT0_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT0_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT0_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT0_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    GT0_RXPCSRESET_IN                       : in   std_logic;
    GT0_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    GT0_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT0_TXUSRCLK_IN                         : in   std_logic;
    GT0_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT0_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT0_GTXTXN_OUT                          : out  std_logic;
    GT0_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT0_TXOUTCLK_OUT                        : out  std_logic;
    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT0_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT0_TXRESETDONE_OUT                     : out  std_logic;

    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT1_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT1_CPLLLOCK_OUT                        : out  std_logic;
    GT1_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT1_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT1_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT1_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT1_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT1_DRPCLK_IN                           : in   std_logic;
    GT1_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT1_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT1_DRPEN_IN                            : in   std_logic;
    GT1_DRPRDY_OUT                          : out  std_logic;
    GT1_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT1_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT1_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT1_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT1_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT1_RXUSRCLK_IN                         : in   std_logic;
    GT1_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT1_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT1_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT1_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT1_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT1_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT1_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT1_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT1_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT1_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT1_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT1_GTRXRESET_IN                        : in   std_logic;
    GT1_RXPCSRESET_IN                       : in   std_logic;
    GT1_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT1_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT1_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT1_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT1_GTTXRESET_IN                        : in   std_logic;
    GT1_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT1_TXUSRCLK_IN                         : in   std_logic;
    GT1_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT1_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT1_GTXTXN_OUT                          : out  std_logic;
    GT1_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT1_TXOUTCLK_OUT                        : out  std_logic;
    GT1_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT1_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT1_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT1_TXRESETDONE_OUT                     : out  std_logic;

    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT2_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT2_CPLLLOCK_OUT                        : out  std_logic;
    GT2_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT2_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT2_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT2_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT2_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT2_DRPCLK_IN                           : in   std_logic;
    GT2_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT2_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT2_DRPEN_IN                            : in   std_logic;
    GT2_DRPRDY_OUT                          : out  std_logic;
    GT2_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT2_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT2_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT2_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT2_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT2_RXUSRCLK_IN                         : in   std_logic;
    GT2_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT2_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT2_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT2_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT2_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT2_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT2_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT2_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT2_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT2_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT2_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT2_GTRXRESET_IN                        : in   std_logic;
    GT2_RXPCSRESET_IN                       : in   std_logic;
    GT2_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT2_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT2_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT2_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT2_GTTXRESET_IN                        : in   std_logic;
    GT2_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT2_TXUSRCLK_IN                         : in   std_logic;
    GT2_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT2_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT2_GTXTXN_OUT                          : out  std_logic;
    GT2_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT2_TXOUTCLK_OUT                        : out  std_logic;
    GT2_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT2_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT2_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT2_TXRESETDONE_OUT                     : out  std_logic;

    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT3_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT3_CPLLLOCK_OUT                        : out  std_logic;
    GT3_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT3_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT3_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT3_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT3_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT3_DRPCLK_IN                           : in   std_logic;
    GT3_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT3_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT3_DRPEN_IN                            : in   std_logic;
    GT3_DRPRDY_OUT                          : out  std_logic;
    GT3_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT3_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT3_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT3_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT3_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT3_RXUSRCLK_IN                         : in   std_logic;
    GT3_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT3_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT3_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT3_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT3_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT3_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT3_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT3_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT3_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT3_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT3_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT3_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT3_GTRXRESET_IN                        : in   std_logic;
    GT3_RXPCSRESET_IN                       : in   std_logic;
    GT3_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT3_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT3_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT3_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT3_GTTXRESET_IN                        : in   std_logic;
    GT3_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT3_TXUSRCLK_IN                         : in   std_logic;
    GT3_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT3_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT3_GTXTXN_OUT                          : out  std_logic;
    GT3_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT3_TXOUTCLK_OUT                        : out  std_logic;
    GT3_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT3_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT3_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT3_TXRESETDONE_OUT                     : out  std_logic;

    --GT4  (X0Y4)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT4_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT4_CPLLLOCK_OUT                        : out  std_logic;
    GT4_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT4_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT4_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT4_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT4_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT4_DRPCLK_IN                           : in   std_logic;
    GT4_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT4_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT4_DRPEN_IN                            : in   std_logic;
    GT4_DRPRDY_OUT                          : out  std_logic;
    GT4_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT4_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT4_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT4_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT4_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT4_RXUSRCLK_IN                         : in   std_logic;
    GT4_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT4_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT4_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT4_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT4_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT4_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT4_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT4_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT4_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT4_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT4_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT4_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT4_GTRXRESET_IN                        : in   std_logic;
    GT4_RXPCSRESET_IN                       : in   std_logic;
    GT4_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT4_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT4_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT4_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT4_GTTXRESET_IN                        : in   std_logic;
    GT4_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT4_TXUSRCLK_IN                         : in   std_logic;
    GT4_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT4_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT4_GTXTXN_OUT                          : out  std_logic;
    GT4_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT4_TXOUTCLK_OUT                        : out  std_logic;
    GT4_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT4_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT4_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT4_TXRESETDONE_OUT                     : out  std_logic;

    --GT5  (X0Y5)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT5_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT5_CPLLLOCK_OUT                        : out  std_logic;
    GT5_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT5_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT5_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT5_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT5_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT5_DRPCLK_IN                           : in   std_logic;
    GT5_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT5_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT5_DRPEN_IN                            : in   std_logic;
    GT5_DRPRDY_OUT                          : out  std_logic;
    GT5_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT5_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT5_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT5_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT5_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT5_RXUSRCLK_IN                         : in   std_logic;
    GT5_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT5_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT5_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT5_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT5_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT5_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT5_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT5_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT5_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT5_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT5_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT5_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT5_GTRXRESET_IN                        : in   std_logic;
    GT5_RXPCSRESET_IN                       : in   std_logic;
    GT5_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT5_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT5_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT5_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT5_GTTXRESET_IN                        : in   std_logic;
    GT5_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT5_TXUSRCLK_IN                         : in   std_logic;
    GT5_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT5_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT5_GTXTXN_OUT                          : out  std_logic;
    GT5_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT5_TXOUTCLK_OUT                        : out  std_logic;
    GT5_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT5_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT5_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT5_TXRESETDONE_OUT                     : out  std_logic;

    --GT6  (X0Y6)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT6_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT6_CPLLLOCK_OUT                        : out  std_logic;
    GT6_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT6_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT6_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT6_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT6_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT6_DRPCLK_IN                           : in   std_logic;
    GT6_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT6_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT6_DRPEN_IN                            : in   std_logic;
    GT6_DRPRDY_OUT                          : out  std_logic;
    GT6_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT6_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT6_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT6_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT6_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT6_RXUSRCLK_IN                         : in   std_logic;
    GT6_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT6_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT6_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT6_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT6_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT6_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT6_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT6_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT6_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT6_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT6_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT6_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT6_GTRXRESET_IN                        : in   std_logic;
    GT6_RXPCSRESET_IN                       : in   std_logic;
    GT6_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT6_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT6_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT6_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT6_GTTXRESET_IN                        : in   std_logic;
    GT6_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT6_TXUSRCLK_IN                         : in   std_logic;
    GT6_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT6_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT6_GTXTXN_OUT                          : out  std_logic;
    GT6_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT6_TXOUTCLK_OUT                        : out  std_logic;
    GT6_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT6_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT6_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT6_TXRESETDONE_OUT                     : out  std_logic;

    --GT7  (X0Y7)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT7_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT7_CPLLLOCK_OUT                        : out  std_logic;
    GT7_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT7_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT7_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT7_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT7_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT7_DRPCLK_IN                           : in   std_logic;
    GT7_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT7_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT7_DRPEN_IN                            : in   std_logic;
    GT7_DRPRDY_OUT                          : out  std_logic;
    GT7_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT7_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT7_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT7_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT7_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT7_RXUSRCLK_IN                         : in   std_logic;
    GT7_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT7_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT7_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT7_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT7_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT7_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT7_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT7_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT7_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT7_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT7_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT7_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT7_GTRXRESET_IN                        : in   std_logic;
    GT7_RXPCSRESET_IN                       : in   std_logic;
    GT7_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT7_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT7_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT7_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT7_GTTXRESET_IN                        : in   std_logic;
    GT7_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT7_TXUSRCLK_IN                         : in   std_logic;
    GT7_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT7_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT7_GTXTXN_OUT                          : out  std_logic;
    GT7_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT7_TXOUTCLK_OUT                        : out  std_logic;
    GT7_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT7_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT7_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT7_TXRESETDONE_OUT                     : out  std_logic;

    --GT8  (X0Y8)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT8_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT8_CPLLLOCK_OUT                        : out  std_logic;
    GT8_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT8_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT8_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT8_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT8_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT8_DRPCLK_IN                           : in   std_logic;
    GT8_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT8_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT8_DRPEN_IN                            : in   std_logic;
    GT8_DRPRDY_OUT                          : out  std_logic;
    GT8_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT8_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT8_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT8_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT8_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT8_RXUSRCLK_IN                         : in   std_logic;
    GT8_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT8_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT8_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT8_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT8_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT8_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT8_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT8_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT8_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT8_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT8_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT8_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT8_GTRXRESET_IN                        : in   std_logic;
    GT8_RXPCSRESET_IN                       : in   std_logic;
    GT8_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT8_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT8_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT8_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT8_GTTXRESET_IN                        : in   std_logic;
    GT8_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT8_TXUSRCLK_IN                         : in   std_logic;
    GT8_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT8_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT8_GTXTXN_OUT                          : out  std_logic;
    GT8_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT8_TXOUTCLK_OUT                        : out  std_logic;
    GT8_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT8_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT8_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT8_TXRESETDONE_OUT                     : out  std_logic;

    --GT9  (X0Y9)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT9_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT9_CPLLLOCK_OUT                        : out  std_logic;
    GT9_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT9_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT9_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT9_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT9_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT9_DRPCLK_IN                           : in   std_logic;
    GT9_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT9_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT9_DRPEN_IN                            : in   std_logic;
    GT9_DRPRDY_OUT                          : out  std_logic;
    GT9_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT9_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT9_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT9_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT9_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT9_RXUSRCLK_IN                         : in   std_logic;
    GT9_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT9_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT9_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT9_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT9_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT9_GTXRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT9_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT9_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT9_RXCOMMADET_OUT                      : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT9_RXDFEAGCHOLD_IN                     : in   std_logic;
    GT9_RXDFELFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT9_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT9_GTRXRESET_IN                        : in   std_logic;
    GT9_RXPCSRESET_IN                       : in   std_logic;
    GT9_RXPMARESET_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT9_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT9_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT9_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT9_GTTXRESET_IN                        : in   std_logic;
    GT9_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT9_TXUSRCLK_IN                         : in   std_logic;
    GT9_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT9_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT9_GTXTXN_OUT                          : out  std_logic;
    GT9_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT9_TXOUTCLK_OUT                        : out  std_logic;
    GT9_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT9_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT9_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT9_TXRESETDONE_OUT                     : out  std_logic;

    --GT10  (X0Y10)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT10_CPLLFBCLKLOST_OUT                  : out  std_logic;
    GT10_CPLLLOCK_OUT                       : out  std_logic;
    GT10_CPLLLOCKDETCLK_IN                  : in   std_logic;
    GT10_CPLLREFCLKLOST_OUT                 : out  std_logic;
    GT10_CPLLRESET_IN                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT10_GTREFCLK0_IN                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT10_DRPADDR_IN                         : in   std_logic_vector(8 downto 0);
    GT10_DRPCLK_IN                          : in   std_logic;
    GT10_DRPDI_IN                           : in   std_logic_vector(15 downto 0);
    GT10_DRPDO_OUT                          : out  std_logic_vector(15 downto 0);
    GT10_DRPEN_IN                           : in   std_logic;
    GT10_DRPRDY_OUT                         : out  std_logic;
    GT10_DRPWE_IN                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT10_LOOPBACK_IN                        : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT10_RXUSERRDY_IN                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT10_EYESCANDATAERROR_OUT               : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT10_RXCDRLOCK_OUT                      : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT10_RXUSRCLK_IN                        : in   std_logic;
    GT10_RXUSRCLK2_IN                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT10_RXDATA_OUT                         : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT10_RXDISPERR_OUT                      : out  std_logic_vector(1 downto 0);
    GT10_RXNOTINTABLE_OUT                   : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT10_GTXRXP_IN                          : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT10_GTXRXN_IN                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT10_RXBYTEISALIGNED_OUT                : out  std_logic;
    GT10_RXBYTEREALIGN_OUT                  : out  std_logic;
    GT10_RXCOMMADET_OUT                     : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT10_RXDFEAGCHOLD_IN                    : in   std_logic;
    GT10_RXDFELFHOLD_IN                     : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT10_RXOUTCLK_OUT                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT10_GTRXRESET_IN                       : in   std_logic;
    GT10_RXPCSRESET_IN                      : in   std_logic;
    GT10_RXPMARESET_IN                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT10_RXCHARISCOMMA_OUT                  : out  std_logic_vector(1 downto 0);
    GT10_RXCHARISK_OUT                      : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT10_RXRESETDONE_OUT                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT10_GTTXRESET_IN                       : in   std_logic;
    GT10_TXUSERRDY_IN                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT10_TXUSRCLK_IN                        : in   std_logic;
    GT10_TXUSRCLK2_IN                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT10_TXDATA_IN                          : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT10_GTXTXN_OUT                         : out  std_logic;
    GT10_GTXTXP_OUT                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT10_TXOUTCLK_OUT                       : out  std_logic;
    GT10_TXOUTCLKFABRIC_OUT                 : out  std_logic;
    GT10_TXOUTCLKPCS_OUT                    : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT10_TXCHARISK_IN                       : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT10_TXRESETDONE_OUT                    : out  std_logic;

    --GT11  (X0Y11)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT11_CPLLFBCLKLOST_OUT                  : out  std_logic;
    GT11_CPLLLOCK_OUT                       : out  std_logic;
    GT11_CPLLLOCKDETCLK_IN                  : in   std_logic;
    GT11_CPLLREFCLKLOST_OUT                 : out  std_logic;
    GT11_CPLLRESET_IN                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT11_GTREFCLK0_IN                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT11_DRPADDR_IN                         : in   std_logic_vector(8 downto 0);
    GT11_DRPCLK_IN                          : in   std_logic;
    GT11_DRPDI_IN                           : in   std_logic_vector(15 downto 0);
    GT11_DRPDO_OUT                          : out  std_logic_vector(15 downto 0);
    GT11_DRPEN_IN                           : in   std_logic;
    GT11_DRPRDY_OUT                         : out  std_logic;
    GT11_DRPWE_IN                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT11_LOOPBACK_IN                        : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT11_RXUSERRDY_IN                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT11_EYESCANDATAERROR_OUT               : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT11_RXCDRLOCK_OUT                      : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT11_RXUSRCLK_IN                        : in   std_logic;
    GT11_RXUSRCLK2_IN                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT11_RXDATA_OUT                         : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT11_RXDISPERR_OUT                      : out  std_logic_vector(1 downto 0);
    GT11_RXNOTINTABLE_OUT                   : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT11_GTXRXP_IN                          : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT11_GTXRXN_IN                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT11_RXBYTEISALIGNED_OUT                : out  std_logic;
    GT11_RXBYTEREALIGN_OUT                  : out  std_logic;
    GT11_RXCOMMADET_OUT                     : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT11_RXDFEAGCHOLD_IN                    : in   std_logic;
    GT11_RXDFELFHOLD_IN                     : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT11_RXOUTCLK_OUT                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT11_GTRXRESET_IN                       : in   std_logic;
    GT11_RXPCSRESET_IN                      : in   std_logic;
    GT11_RXPMARESET_IN                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT11_RXCHARISCOMMA_OUT                  : out  std_logic_vector(1 downto 0);
    GT11_RXCHARISK_OUT                      : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT11_RXRESETDONE_OUT                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT11_GTTXRESET_IN                       : in   std_logic;
    GT11_TXUSERRDY_IN                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT11_TXUSRCLK_IN                        : in   std_logic;
    GT11_TXUSRCLK2_IN                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT11_TXDATA_IN                          : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT11_GTXTXN_OUT                         : out  std_logic;
    GT11_GTXTXP_OUT                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT11_TXOUTCLK_OUT                       : out  std_logic;
    GT11_TXOUTCLKFABRIC_OUT                 : out  std_logic;
    GT11_TXOUTCLKPCS_OUT                    : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT11_TXCHARISK_IN                       : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT11_TXRESETDONE_OUT                    : out  std_logic;


    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    GT0_GTREFCLK0_COMMON_IN                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    GT0_QPLLLOCK_OUT                        : out  std_logic;
    GT0_QPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_QPLLREFCLKLOST_OUT                  : out  std_logic;
    GT0_QPLLRESET_IN                        : in   std_logic;

    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    GT1_GTREFCLK0_COMMON_IN                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    GT1_QPLLLOCK_OUT                        : out  std_logic;
    GT1_QPLLLOCKDETCLK_IN                   : in   std_logic;
    GT1_QPLLREFCLKLOST_OUT                  : out  std_logic;
    GT1_QPLLRESET_IN                        : in   std_logic;

    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    GT2_GTREFCLK0_COMMON_IN                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    GT2_QPLLLOCK_OUT                        : out  std_logic;
    GT2_QPLLLOCKDETCLK_IN                   : in   std_logic;
    GT2_QPLLREFCLKLOST_OUT                  : out  std_logic;
    GT2_QPLLRESET_IN                        : in   std_logic


);


end gtx_minipod_12x_k7;
    
architecture RTL of gtx_minipod_12x_k7 is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gtx_minipod_12x_k7,gtwizard_v2_6,{protocol_file=Start_from_scratch}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;
    signal   gt0_qplloutclk_i         :   std_logic;
    signal   gt0_qplloutrefclk_i      :   std_logic;
    signal   gt1_qplloutclk_i         :   std_logic;
    signal   gt1_qplloutrefclk_i      :   std_logic;
    signal   gt2_qplloutclk_i         :   std_logic;
    signal   gt2_qplloutrefclk_i      :   std_logic;

  
    signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt4_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt4_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt5_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt5_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt6_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt6_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt7_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt7_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt8_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt8_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt9_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt9_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt10_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt10_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt11_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt11_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
 
    signal   gt0_qpllclk_i            :   std_logic;
    signal   gt0_qpllrefclk_i         :   std_logic;
    signal   gt1_qpllclk_i            :   std_logic;
    signal   gt1_qpllrefclk_i         :   std_logic;
    signal   gt2_qpllclk_i            :   std_logic;
    signal   gt2_qpllrefclk_i         :   std_logic;
    signal   gt3_qpllclk_i            :   std_logic;
    signal   gt3_qpllrefclk_i         :   std_logic;
    signal   gt4_qpllclk_i            :   std_logic;
    signal   gt4_qpllrefclk_i         :   std_logic;
    signal   gt5_qpllclk_i            :   std_logic;
    signal   gt5_qpllrefclk_i         :   std_logic;
    signal   gt6_qpllclk_i            :   std_logic;
    signal   gt6_qpllrefclk_i         :   std_logic;
    signal   gt7_qpllclk_i            :   std_logic;
    signal   gt7_qpllrefclk_i         :   std_logic;
    signal   gt8_qpllclk_i            :   std_logic;
    signal   gt8_qpllrefclk_i         :   std_logic;
    signal   gt9_qpllclk_i            :   std_logic;
    signal   gt9_qpllrefclk_i         :   std_logic;
    signal   gt10_qpllclk_i            :   std_logic;
    signal   gt10_qpllrefclk_i         :   std_logic;
    signal   gt11_qpllclk_i            :   std_logic;
    signal   gt11_qpllrefclk_i         :   std_logic;


--*************************** Component Declarations **************************
component gtx_minipod_12x_k7_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP       : string   := "FALSE";
    RX_DFE_KL_CFG2_IN            : bit_vector :=   X"3010D90C";
    PMA_RSV_IN                   : bit_vector :=   X"00000000";
    PCS_RSVD_ATTR_IN             : bit_vector :=   X"000000000000"
);
port 
(   
    --------------------------------- CPLL Ports -------------------------------
    CPLLFBCLKLOST_OUT                       : out  std_logic;
    CPLLLOCK_OUT                            : out  std_logic;
    CPLLLOCKDETCLK_IN                       : in   std_logic;
    CPLLREFCLKLOST_OUT                      : out  std_logic;
    CPLLRESET_IN                            : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GTREFCLK0_IN                            : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    DRPADDR_IN                              : in   std_logic_vector(8 downto 0);
    DRPCLK_IN                               : in   std_logic;
    DRPDI_IN                                : in   std_logic_vector(15 downto 0);
    DRPDO_OUT                               : out  std_logic_vector(15 downto 0);
    DRPEN_IN                                : in   std_logic;
    DRPRDY_OUT                              : out  std_logic;
    DRPWE_IN                                : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    QPLLCLK_IN                              : in   std_logic;
    QPLLREFCLK_IN                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    LOOPBACK_IN                             : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    RXUSERRDY_IN                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    EYESCANDATAERROR_OUT                    : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    RXCDRLOCK_OUT                           : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    RXUSRCLK_IN                             : in   std_logic;
    RXUSRCLK2_IN                            : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    RXDATA_OUT                              : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    RXDISPERR_OUT                           : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE_OUT                        : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GTXRXP_IN                               : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GTXRXN_IN                               : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    RXBYTEISALIGNED_OUT                     : out  std_logic;
    RXBYTEREALIGN_OUT                       : out  std_logic;
    RXCOMMADET_OUT                          : out  std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    RXDFEAGCHOLD_IN                         : in   std_logic;
    RXDFELFHOLD_IN                          : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    RXOUTCLK_OUT                            : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GTRXRESET_IN                            : in   std_logic;
    RXPCSRESET_IN                           : in   std_logic;
    RXPMARESET_IN                           : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    RXCHARISCOMMA_OUT                       : out  std_logic_vector(1 downto 0);
    RXCHARISK_OUT                           : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    RXRESETDONE_OUT                         : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GTTXRESET_IN                            : in   std_logic;
    TXUSERRDY_IN                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    TXUSRCLK_IN                             : in   std_logic;
    TXUSRCLK2_IN                            : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TXDATA_IN                               : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTXTXN_OUT                              : out  std_logic;
    GTXTXP_OUT                              : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    TXOUTCLK_OUT                            : out  std_logic;
    TXOUTCLKFABRIC_OUT                      : out  std_logic;
    TXOUTCLKPCS_OUT                         : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    TXCHARISK_IN                            : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    TXRESETDONE_OUT                         : out  std_logic


);
end component;



--*************************Logic to set Attribute QPLL_FB_DIV*****************************
    impure function conv_qpll_fbdiv_top (qpllfbdiv_top : in integer) return bit_vector is
    begin
       if (qpllfbdiv_top = 16) then
         return "0000100000";
       elsif (qpllfbdiv_top = 20) then
         return "0000110000" ;
       elsif (qpllfbdiv_top = 32) then
         return "0001100000" ;
       elsif (qpllfbdiv_top = 40) then
         return "0010000000" ;
       elsif (qpllfbdiv_top = 64) then
         return "0011100000" ;
       elsif (qpllfbdiv_top = 66) then
         return "0101000000" ;
       elsif (qpllfbdiv_top = 80) then
         return "0100100000" ;
       elsif (qpllfbdiv_top = 100) then
         return "0101110000" ;
       else 
         return "0000000000" ;
       end if;
    end function;

    impure function conv_qpll_fbdiv_ratio (qpllfbdiv_top : in integer) return bit is
    begin
       if (qpllfbdiv_top = 16) then
         return '1';
       elsif (qpllfbdiv_top = 20) then
         return '1' ;
       elsif (qpllfbdiv_top = 32) then
         return '1' ;
       elsif (qpllfbdiv_top = 40) then
         return '1' ;
       elsif (qpllfbdiv_top = 64) then
         return '1' ;
       elsif (qpllfbdiv_top = 66) then
         return '0' ;
       elsif (qpllfbdiv_top = 80) then
         return '1' ;
       elsif (qpllfbdiv_top = 100) then
         return '1' ;
       else 
         return '1' ;
       end if;
    end function;

    constant   QPLL_FBDIV_IN    :   bit_vector(9 downto 0) := conv_qpll_fbdiv_top(QPLL_FBDIV_TOP);
    constant   QPLL_FBDIV_RATIO :   bit := conv_qpll_fbdiv_ratio(QPLL_FBDIV_TOP);

--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_qpllclk_i    <= gt0_qplloutclk_i;  
    gt0_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt1_qpllclk_i    <= gt0_qplloutclk_i;  
    gt1_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt2_qpllclk_i    <= gt0_qplloutclk_i;  
    gt2_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt3_qpllclk_i    <= gt0_qplloutclk_i;  
    gt3_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt4_qpllclk_i    <= gt1_qplloutclk_i;  
    gt4_qpllrefclk_i <= gt1_qplloutrefclk_i; 

    gt5_qpllclk_i    <= gt1_qplloutclk_i;  
    gt5_qpllrefclk_i <= gt1_qplloutrefclk_i; 

    gt6_qpllclk_i    <= gt1_qplloutclk_i;  
    gt6_qpllrefclk_i <= gt1_qplloutrefclk_i; 

    gt7_qpllclk_i    <= gt1_qplloutclk_i;  
    gt7_qpllrefclk_i <= gt1_qplloutrefclk_i; 

    gt8_qpllclk_i    <= gt2_qplloutclk_i;  
    gt8_qpllrefclk_i <= gt2_qplloutrefclk_i; 

    gt9_qpllclk_i    <= gt2_qplloutclk_i;  
    gt9_qpllrefclk_i <= gt2_qplloutrefclk_i; 

    gt10_qpllclk_i    <= gt2_qplloutclk_i;  
    gt10_qpllrefclk_i <= gt2_qplloutrefclk_i; 

    gt11_qpllclk_i    <= gt2_qplloutclk_i;  
    gt11_qpllrefclk_i <= gt2_qplloutrefclk_i; 


 
    --------------------------- GT Instances  -------------------------------   

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)

    gt0_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT0_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT0_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT0_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT0_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT0_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT0_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT0_DRPADDR_IN,
        DRPCLK_IN                       =>      GT0_DRPCLK_IN,
        DRPDI_IN                        =>      GT0_DRPDI_IN,
        DRPDO_OUT                       =>      GT0_DRPDO_OUT,
        DRPEN_IN                        =>      GT0_DRPEN_IN,
        DRPRDY_OUT                      =>      GT0_DRPRDY_OUT,
        DRPWE_IN                        =>      GT0_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt0_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt0_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT0_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT0_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT0_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT0_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT0_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT0_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT0_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT0_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT0_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT0_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT0_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT0_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT0_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT0_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT0_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT0_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT0_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT0_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT0_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT0_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT0_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT0_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT0_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT0_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT0_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT0_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT0_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT0_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT0_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT0_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT0_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT0_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT0_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT0_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT0_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y1)

    gt1_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT1_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT1_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT1_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT1_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT1_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT1_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT1_DRPADDR_IN,
        DRPCLK_IN                       =>      GT1_DRPCLK_IN,
        DRPDI_IN                        =>      GT1_DRPDI_IN,
        DRPDO_OUT                       =>      GT1_DRPDO_OUT,
        DRPEN_IN                        =>      GT1_DRPEN_IN,
        DRPRDY_OUT                      =>      GT1_DRPRDY_OUT,
        DRPWE_IN                        =>      GT1_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt1_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt1_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT1_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT1_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT1_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT1_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT1_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT1_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT1_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT1_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT1_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT1_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT1_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT1_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT1_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT1_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT1_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT1_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT1_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT1_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT1_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT1_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT1_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT1_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT1_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT1_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT1_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT1_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT1_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT1_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT1_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT1_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT1_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT1_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT1_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT1_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT1_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y2)

    gt2_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT2_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT2_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT2_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT2_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT2_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT2_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT2_DRPADDR_IN,
        DRPCLK_IN                       =>      GT2_DRPCLK_IN,
        DRPDI_IN                        =>      GT2_DRPDI_IN,
        DRPDO_OUT                       =>      GT2_DRPDO_OUT,
        DRPEN_IN                        =>      GT2_DRPEN_IN,
        DRPRDY_OUT                      =>      GT2_DRPRDY_OUT,
        DRPWE_IN                        =>      GT2_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt2_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt2_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT2_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT2_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT2_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT2_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT2_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT2_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT2_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT2_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT2_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT2_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT2_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT2_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT2_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT2_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT2_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT2_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT2_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT2_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT2_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT2_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT2_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT2_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT2_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT2_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT2_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT2_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT2_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT2_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT2_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT2_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT2_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT2_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT2_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT2_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT2_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y3)

    gt3_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT3_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT3_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT3_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT3_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT3_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT3_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT3_DRPADDR_IN,
        DRPCLK_IN                       =>      GT3_DRPCLK_IN,
        DRPDI_IN                        =>      GT3_DRPDI_IN,
        DRPDO_OUT                       =>      GT3_DRPDO_OUT,
        DRPEN_IN                        =>      GT3_DRPEN_IN,
        DRPRDY_OUT                      =>      GT3_DRPRDY_OUT,
        DRPWE_IN                        =>      GT3_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt3_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt3_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT3_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT3_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT3_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT3_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT3_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT3_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT3_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT3_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT3_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT3_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT3_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT3_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT3_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT3_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT3_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT3_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT3_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT3_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT3_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT3_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT3_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT3_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT3_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT3_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT3_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT3_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT3_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT3_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT3_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT3_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT3_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT3_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT3_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT3_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT3_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT4  (X0Y4)

    gt4_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT4_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT4_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT4_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT4_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT4_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT4_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT4_DRPADDR_IN,
        DRPCLK_IN                       =>      GT4_DRPCLK_IN,
        DRPDI_IN                        =>      GT4_DRPDI_IN,
        DRPDO_OUT                       =>      GT4_DRPDO_OUT,
        DRPEN_IN                        =>      GT4_DRPEN_IN,
        DRPRDY_OUT                      =>      GT4_DRPRDY_OUT,
        DRPWE_IN                        =>      GT4_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt4_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt4_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT4_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT4_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT4_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT4_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT4_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT4_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT4_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT4_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT4_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT4_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT4_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT4_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT4_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT4_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT4_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT4_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT4_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT4_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT4_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT4_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT4_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT4_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT4_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT4_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT4_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT4_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT4_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT4_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT4_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT4_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT4_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT4_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT4_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT4_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT4_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT5  (X0Y5)

    gt5_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT5_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT5_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT5_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT5_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT5_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT5_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT5_DRPADDR_IN,
        DRPCLK_IN                       =>      GT5_DRPCLK_IN,
        DRPDI_IN                        =>      GT5_DRPDI_IN,
        DRPDO_OUT                       =>      GT5_DRPDO_OUT,
        DRPEN_IN                        =>      GT5_DRPEN_IN,
        DRPRDY_OUT                      =>      GT5_DRPRDY_OUT,
        DRPWE_IN                        =>      GT5_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt5_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt5_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT5_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT5_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT5_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT5_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT5_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT5_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT5_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT5_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT5_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT5_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT5_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT5_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT5_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT5_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT5_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT5_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT5_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT5_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT5_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT5_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT5_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT5_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT5_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT5_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT5_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT5_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT5_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT5_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT5_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT5_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT5_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT5_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT5_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT5_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT5_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT6  (X0Y6)

    gt6_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT6_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT6_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT6_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT6_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT6_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT6_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT6_DRPADDR_IN,
        DRPCLK_IN                       =>      GT6_DRPCLK_IN,
        DRPDI_IN                        =>      GT6_DRPDI_IN,
        DRPDO_OUT                       =>      GT6_DRPDO_OUT,
        DRPEN_IN                        =>      GT6_DRPEN_IN,
        DRPRDY_OUT                      =>      GT6_DRPRDY_OUT,
        DRPWE_IN                        =>      GT6_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt6_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt6_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT6_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT6_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT6_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT6_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT6_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT6_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT6_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT6_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT6_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT6_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT6_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT6_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT6_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT6_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT6_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT6_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT6_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT6_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT6_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT6_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT6_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT6_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT6_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT6_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT6_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT6_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT6_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT6_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT6_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT6_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT6_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT6_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT6_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT6_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT6_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT7  (X0Y7)

    gt7_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT7_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT7_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT7_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT7_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT7_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT7_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT7_DRPADDR_IN,
        DRPCLK_IN                       =>      GT7_DRPCLK_IN,
        DRPDI_IN                        =>      GT7_DRPDI_IN,
        DRPDO_OUT                       =>      GT7_DRPDO_OUT,
        DRPEN_IN                        =>      GT7_DRPEN_IN,
        DRPRDY_OUT                      =>      GT7_DRPRDY_OUT,
        DRPWE_IN                        =>      GT7_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt7_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt7_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT7_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT7_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT7_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT7_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT7_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT7_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT7_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT7_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT7_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT7_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT7_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT7_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT7_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT7_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT7_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT7_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT7_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT7_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT7_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT7_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT7_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT7_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT7_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT7_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT7_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT7_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT7_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT7_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT7_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT7_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT7_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT7_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT7_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT7_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT7_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT8  (X0Y8)

    gt8_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT8_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT8_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT8_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT8_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT8_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT8_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT8_DRPADDR_IN,
        DRPCLK_IN                       =>      GT8_DRPCLK_IN,
        DRPDI_IN                        =>      GT8_DRPDI_IN,
        DRPDO_OUT                       =>      GT8_DRPDO_OUT,
        DRPEN_IN                        =>      GT8_DRPEN_IN,
        DRPRDY_OUT                      =>      GT8_DRPRDY_OUT,
        DRPWE_IN                        =>      GT8_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt8_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt8_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT8_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT8_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT8_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT8_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT8_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT8_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT8_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT8_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT8_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT8_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT8_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT8_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT8_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT8_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT8_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT8_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT8_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT8_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT8_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT8_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT8_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT8_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT8_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT8_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT8_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT8_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT8_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT8_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT8_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT8_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT8_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT8_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT8_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT8_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT8_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT9  (X0Y9)

    gt9_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT9_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT9_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT9_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT9_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT9_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT9_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT9_DRPADDR_IN,
        DRPCLK_IN                       =>      GT9_DRPCLK_IN,
        DRPDI_IN                        =>      GT9_DRPDI_IN,
        DRPDO_OUT                       =>      GT9_DRPDO_OUT,
        DRPEN_IN                        =>      GT9_DRPEN_IN,
        DRPRDY_OUT                      =>      GT9_DRPRDY_OUT,
        DRPWE_IN                        =>      GT9_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt9_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt9_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT9_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT9_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT9_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT9_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT9_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT9_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT9_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT9_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT9_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT9_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT9_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT9_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT9_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT9_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT9_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT9_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT9_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT9_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT9_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT9_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT9_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT9_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT9_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT9_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT9_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT9_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT9_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT9_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT9_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT9_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT9_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT9_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT9_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT9_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT9_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT10  (X0Y10)

    gt10_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT10_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT10_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT10_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT10_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT10_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT10_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT10_DRPADDR_IN,
        DRPCLK_IN                       =>      GT10_DRPCLK_IN,
        DRPDI_IN                        =>      GT10_DRPDI_IN,
        DRPDO_OUT                       =>      GT10_DRPDO_OUT,
        DRPEN_IN                        =>      GT10_DRPEN_IN,
        DRPRDY_OUT                      =>      GT10_DRPRDY_OUT,
        DRPWE_IN                        =>      GT10_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt10_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt10_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT10_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT10_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT10_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT10_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT10_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT10_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT10_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT10_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT10_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT10_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT10_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT10_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT10_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT10_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT10_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT10_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT10_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT10_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT10_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT10_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT10_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT10_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT10_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT10_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT10_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT10_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT10_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT10_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT10_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT10_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT10_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT10_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT10_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT10_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT10_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT11  (X0Y11)

    gt11_gtx_minipod_12x_k7_i : gtx_minipod_12x_k7_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000"
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT11_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT11_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT11_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT11_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT11_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT11_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT11_DRPADDR_IN,
        DRPCLK_IN                       =>      GT11_DRPCLK_IN,
        DRPDI_IN                        =>      GT11_DRPDI_IN,
        DRPDO_OUT                       =>      GT11_DRPDO_OUT,
        DRPEN_IN                        =>      GT11_DRPEN_IN,
        DRPRDY_OUT                      =>      GT11_DRPRDY_OUT,
        DRPWE_IN                        =>      GT11_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt11_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt11_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        LOOPBACK_IN                     =>      GT11_LOOPBACK_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT11_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT11_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRLOCK_OUT                   =>      GT11_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT11_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT11_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT11_RXDATA_OUT,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        RXDISPERR_OUT                   =>      GT11_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT11_RXNOTINTABLE_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT11_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT11_GTXRXN_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        RXBYTEISALIGNED_OUT             =>      GT11_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT11_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT11_RXCOMMADET_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFEAGCHOLD_IN                 =>      GT11_RXDFEAGCHOLD_IN,
        RXDFELFHOLD_IN                  =>      GT11_RXDFELFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT11_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT11_GTRXRESET_IN,
        RXPCSRESET_IN                   =>      GT11_RXPCSRESET_IN,
        RXPMARESET_IN                   =>      GT11_RXPMARESET_IN,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        RXCHARISCOMMA_OUT               =>      GT11_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT11_RXCHARISK_OUT,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT11_RXRESETDONE_OUT,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT11_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT11_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT11_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT11_TXUSRCLK2_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT11_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT11_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT11_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT11_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT11_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT11_TXOUTCLKPCS_OUT,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        TXCHARISK_IN                    =>      GT11_TXCHARISK_IN,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXRESETDONE_OUT                 =>      GT11_TXRESETDONE_OUT

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --_________________________GTXE2_COMMON____________________________________

    gtxe2_common_0_i : GTXE2_COMMON
    generic map
    (
            -- Simulation attributes
            SIM_RESET_SPEEDUP    => WRAPPER_SIM_GTRESET_SPEEDUP,
            SIM_QPLLREFCLK_SEL   => ("001"),
            SIM_VERSION          => "4.0",


       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000040000001000"),
        COMMON_CFG                              =>     (x"00000000"),
        QPLL_CFG                                =>     (x"06801C1"),
        QPLL_CLKOUT_CFG                         =>     ("0000"),
        QPLL_COARSE_FREQ_OVRD                   =>     ("010000"),
        QPLL_COARSE_FREQ_OVRD_EN                =>     ('0'),
        QPLL_CP                                 =>     ("0000011111"),
        QPLL_CP_MONITOR_EN                      =>     ('0'),
        QPLL_DMONITOR_SEL                       =>     ('0'),
        QPLL_FBDIV                              =>     (QPLL_FBDIV_IN),
        QPLL_FBDIV_MONITOR_EN                   =>     ('0'),
        QPLL_FBDIV_RATIO                        =>     (QPLL_FBDIV_RATIO),
        QPLL_INIT_CFG                           =>     (x"000006"),
        QPLL_LOCK_CFG                           =>     (x"21E8"),
        QPLL_LPF                                =>     ("1111"),
        QPLL_REFCLK_DIV                         =>     (1)

        
    )
    port map
    (
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GTGREFCLK                       =>      tied_to_ground_i,
        GTNORTHREFCLK0                  =>      tied_to_ground_i,
        GTNORTHREFCLK1                  =>      tied_to_ground_i,
        GTREFCLK0                       =>      GT0_GTREFCLK0_COMMON_IN,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTSOUTHREFCLK0                  =>      tied_to_ground_i,
        GTSOUTHREFCLK1                  =>      tied_to_ground_i,
        ------------------------- Common Block -  QPLL Ports -----------------------
        QPLLDMONITOR                    =>      open,
        ----------------------- Common Block - Clocking Ports ----------------------
        QPLLOUTCLK                      =>      gt0_qplloutclk_i,
        QPLLOUTREFCLK                   =>      gt0_qplloutrefclk_i,
        REFCLKOUTMONITOR                =>      open,
        ------------------------- Common Block - QPLL Ports ------------------------
        QPLLFBCLKLOST                   =>      open,
        QPLLLOCK                        =>      GT0_QPLLLOCK_OUT,
        QPLLLOCKDETCLK                  =>      GT0_QPLLLOCKDETCLK_IN,
        QPLLLOCKEN                      =>      tied_to_vcc_i,
        QPLLOUTRESET                    =>      tied_to_ground_i,
        QPLLPD                          =>      tied_to_ground_i,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_OUT,
        QPLLREFCLKSEL                   =>      "001",
        QPLLRESET                       =>      GT0_QPLLRESET_IN,
        QPLLRSVD1                       =>      "0000000000000000",
        QPLLRSVD2                       =>      "11111",
        --------------------------------- QPLL Ports -------------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i

    );


    --_________________________________________________________________________
    --_________________________________________________________________________
    --_________________________GTXE2_COMMON____________________________________

    gtxe2_common_1_i : GTXE2_COMMON
    generic map
    (
            -- Simulation attributes
            SIM_RESET_SPEEDUP    => WRAPPER_SIM_GTRESET_SPEEDUP,
            SIM_QPLLREFCLK_SEL   => ("001"),
            SIM_VERSION          => "4.0",


       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000040000001000"),
        COMMON_CFG                              =>     (x"00000000"),
        QPLL_CFG                                =>     (x"06801C1"),
        QPLL_CLKOUT_CFG                         =>     ("0000"),
        QPLL_COARSE_FREQ_OVRD                   =>     ("010000"),
        QPLL_COARSE_FREQ_OVRD_EN                =>     ('0'),
        QPLL_CP                                 =>     ("0000011111"),
        QPLL_CP_MONITOR_EN                      =>     ('0'),
        QPLL_DMONITOR_SEL                       =>     ('0'),
        QPLL_FBDIV                              =>     (QPLL_FBDIV_IN),
        QPLL_FBDIV_MONITOR_EN                   =>     ('0'),
        QPLL_FBDIV_RATIO                        =>     (QPLL_FBDIV_RATIO),
        QPLL_INIT_CFG                           =>     (x"000006"),
        QPLL_LOCK_CFG                           =>     (x"21E8"),
        QPLL_LPF                                =>     ("1111"),
        QPLL_REFCLK_DIV                         =>     (1)

        
    )
    port map
    (
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GTGREFCLK                       =>      tied_to_ground_i,
        GTNORTHREFCLK0                  =>      tied_to_ground_i,
        GTNORTHREFCLK1                  =>      tied_to_ground_i,
        GTREFCLK0                       =>      GT1_GTREFCLK0_COMMON_IN,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTSOUTHREFCLK0                  =>      tied_to_ground_i,
        GTSOUTHREFCLK1                  =>      tied_to_ground_i,
        ------------------------- Common Block -  QPLL Ports -----------------------
        QPLLDMONITOR                    =>      open,
        ----------------------- Common Block - Clocking Ports ----------------------
        QPLLOUTCLK                      =>      gt1_qplloutclk_i,
        QPLLOUTREFCLK                   =>      gt1_qplloutrefclk_i,
        REFCLKOUTMONITOR                =>      open,
        ------------------------- Common Block - QPLL Ports ------------------------
        QPLLFBCLKLOST                   =>      open,
        QPLLLOCK                        =>      GT1_QPLLLOCK_OUT,
        QPLLLOCKDETCLK                  =>      GT1_QPLLLOCKDETCLK_IN,
        QPLLLOCKEN                      =>      tied_to_vcc_i,
        QPLLOUTRESET                    =>      tied_to_ground_i,
        QPLLPD                          =>      tied_to_ground_i,
        QPLLREFCLKLOST                  =>      GT1_QPLLREFCLKLOST_OUT,
        QPLLREFCLKSEL                   =>      "001",
        QPLLRESET                       =>      GT1_QPLLRESET_IN,
        QPLLRSVD1                       =>      "0000000000000000",
        QPLLRSVD2                       =>      "11111",
        --------------------------------- QPLL Ports -------------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i

    );


    --_________________________________________________________________________
    --_________________________________________________________________________
    --_________________________GTXE2_COMMON____________________________________

    gtxe2_common_2_i : GTXE2_COMMON
    generic map
    (
            -- Simulation attributes
            SIM_RESET_SPEEDUP    => WRAPPER_SIM_GTRESET_SPEEDUP,
            SIM_QPLLREFCLK_SEL   => ("001"),
            SIM_VERSION          => "4.0",


       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000040000001000"),
        COMMON_CFG                              =>     (x"00000000"),
        QPLL_CFG                                =>     (x"06801C1"),
        QPLL_CLKOUT_CFG                         =>     ("0000"),
        QPLL_COARSE_FREQ_OVRD                   =>     ("010000"),
        QPLL_COARSE_FREQ_OVRD_EN                =>     ('0'),
        QPLL_CP                                 =>     ("0000011111"),
        QPLL_CP_MONITOR_EN                      =>     ('0'),
        QPLL_DMONITOR_SEL                       =>     ('0'),
        QPLL_FBDIV                              =>     (QPLL_FBDIV_IN),
        QPLL_FBDIV_MONITOR_EN                   =>     ('0'),
        QPLL_FBDIV_RATIO                        =>     (QPLL_FBDIV_RATIO),
        QPLL_INIT_CFG                           =>     (x"000006"),
        QPLL_LOCK_CFG                           =>     (x"21E8"),
        QPLL_LPF                                =>     ("1111"),
        QPLL_REFCLK_DIV                         =>     (1)

        
    )
    port map
    (
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GTGREFCLK                       =>      tied_to_ground_i,
        GTNORTHREFCLK0                  =>      tied_to_ground_i,
        GTNORTHREFCLK1                  =>      tied_to_ground_i,
        GTREFCLK0                       =>      GT2_GTREFCLK0_COMMON_IN,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTSOUTHREFCLK0                  =>      tied_to_ground_i,
        GTSOUTHREFCLK1                  =>      tied_to_ground_i,
        ------------------------- Common Block -  QPLL Ports -----------------------
        QPLLDMONITOR                    =>      open,
        ----------------------- Common Block - Clocking Ports ----------------------
        QPLLOUTCLK                      =>      gt2_qplloutclk_i,
        QPLLOUTREFCLK                   =>      gt2_qplloutrefclk_i,
        REFCLKOUTMONITOR                =>      open,
        ------------------------- Common Block - QPLL Ports ------------------------
        QPLLFBCLKLOST                   =>      open,
        QPLLLOCK                        =>      GT2_QPLLLOCK_OUT,
        QPLLLOCKDETCLK                  =>      GT2_QPLLLOCKDETCLK_IN,
        QPLLLOCKEN                      =>      tied_to_vcc_i,
        QPLLOUTRESET                    =>      tied_to_ground_i,
        QPLLPD                          =>      tied_to_ground_i,
        QPLLREFCLKLOST                  =>      GT2_QPLLREFCLKLOST_OUT,
        QPLLREFCLKSEL                   =>      "001",
        QPLLRESET                       =>      GT2_QPLLRESET_IN,
        QPLLRSVD1                       =>      "0000000000000000",
        QPLLRSVD2                       =>      "11111",
        --------------------------------- QPLL Ports -------------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i

    );


     
end RTL;
