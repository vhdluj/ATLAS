`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Bap7yrVl+ScwAs+FKOj9pduUFoJ1DQp0mZakC7cmADqm+EV3/AvrcU8oTYjyziFwk0aAKdjkbojL
CZUjZlNnhw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cJrJC1YhUiRkkcz37hx/zr3sNWhiMjg/guM9xpcXOyN8ZhA9f/+GPAf0fk9aKBzTrOd9ojqXxRch
kcpjPoUI/f08TBz7zlhGegb76wMooraLh6sJVFNW09LT4VDgv/6dfNk9i/CJZ4QgyJfEa2F/E1ky
oXiO/iWXU4UAIW73ZRA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
56cXOoSlLVLHiRVaoWF5E16U5FH6Lpe/8aKgIJJ0jeWqMPxsA92492EmPxqSjIFbtsO1TaFYOPSk
lX7u/vXtX6twpeQiGXXo5me+rC4zCmoxZV8AZumNT/JcRx+tcxaZ6lfA3c26AKirfqK20VNjokco
zWeZbz8qbG3hCH6106vrlCbEGDSvERLT1cs8a1ZNGN0tHkIZAoqgUbR7SC2+RvZVW8rqb3zVvr6F
0B4aQ8u1xyxcT1dHxfAHIjdW0ZFJwPaYQqPJ7BIk9KK3Vo7n55ZxkET4Rj/ren4mED2I6SRuyITn
hv+j0aBNvnZWlUoAwwfG5nlUsdqJqox6maYVlg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pCd0hFVzDSlFCf3du9EpSHQOW8CksqXVQGZNHZO3l/wiaWC5L1x4kGvRAoMG9gCdooqG2laxUPUE
sIOrLm4FwBoE8vY0tXEr8UJqYhriOt5PE8pVkIYDTajJlphe51IafDSyzHyAqoQWYYcYVWwaihxH
D7CY12p+WpjaVm548xo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GwiMJF8w0QuK1hx1itQZ7o1zVbo4St6szK0uw2PeUgv6krJXxaJZbCwxGAty1XgqZwtc8nmEa0NE
wvQ6M8fEqm36puJELtr6C6hoSBwnVSnYKS/AEDeN0VDgmHPoBzU1TH2Awumv++pdW/I3o8oeiwGn
lpyMLdnDucIiKAvc1A7a9qJ5gFhEOLNHNswrQPg8AkIpGeEgPi4ASeoH981KAtGgO4SVtADJlkgT
io2S+iz7lSqAjqEG5StfAOzDhNTTWekrNqGiderJE/Y+4H6FvUmc+/5G46To9PUQqnMKW9DAARxq
uC6/5rQ6U0/XQQ0oiDUdtSfKyGbZdtAZMF5k8g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16592)
`protect data_block
m83KgzB+plw0S+OiSBj3NMJbpyMZ0RlVitsB00R0tUGB37lxZg3fnEzGyvfJTRIZa2Hm1Oy7hTDf
o3CJxHwQQxd9f4wRVIRUCoOGz2NMGCxyESMJTVDLjZftKMvwCYEj7R2qx16+VsVs0xN5dAoR4iGn
CE94gZ+KWxrzX33NExCN1ikLbAgOaZEbIMroQaGexKD+KUfyuWg2JAia2wBIsPM88j7jz0oqTH5s
LonQ9Jz4pKEdOhO8VvGNL3lyTewk1rWVga+v0/UP2w99AIykkw93I7HkmDVsaKZGREnDx6NFJ9lr
0YDA0OTPQ5iDuaZ08TlUQ7UbIRkkUFpOVxI+3VMsUacaYMc4H+MCC3R+0GrsJTUQh5cV4gQ0qY+l
EE6wt+uf5Zj8DKpPFG6UiswhyTaTzLQJqfPDKGwp+pggOS3FZXFIsogCqoob7/EFJo6clfMyZWOs
jH5wQxYuffXi+X9rKeJkOphkl2WxUbtyfvdHkx0g8loxqTSYUHpbVnp7Lj2eqDRFJqcEp6svWiNe
f6RKdYx8GFfuuE2PbJDyTjWCCi1yBt53pXYCXnquZHGdSniyhKaKx/G7Mw3lFLzBKqcjT3wsvQtI
dnDFaXzj5C3637KFS6lteT3Bog90YO7pDJXKIuWfyT+nNipieIOkCb1PLbFCmNA895KW8mvF48Cz
hIwfj3AHNXKsE9RKLWiEYS7PGxzYoQ+hx6GfbbMWqLITpqOArK7hjwndoJUvIl+TWSP6rSFsrTOu
JlIPZvBhKSTaUjP8Cjk9D5XFpBrxiqQgcaBPbr4Eg+1fkNMzQwMzecdZpqKy15unowZ9IEkFML+C
bHBJIElICvU5Zsv8JNibjzyNygFqzTlQS3ggRNpU3DmD6TROq9nMhbCcb074dQMevFeS3Dcz0hCj
gTbSMUkWlisrfKnfYN2tOD5jahglzS4efKO1naW5dLZnf6FilrGK2KvHYUa+DKinkMJhJxD7K0Wg
4QFUy4Mw875v+rjjeePD4SMijONHBruzg7yWhryDZrhwlMnwm8coWi2JIMUM/4YLWKBR3Mlrobek
By9dWaJIAXYx9h/uqtwdSgnryX3ZMF7DqzFE2+q1R80w2+/ihd1gSvEjCbB5nZ9SrjeMIlLgfWJP
gYvj8x7YTkQqUq0gVrUqJBcHa9RFgz4KoJeGQuWWBh3HAhLcLslXtot2pzN+xr47enS5gt+DAA18
EJsXMQ9a+1AO1nvKHvUMblhZZb1YuVzExmocX+D1hiomuDG3QGOg93h63QkT8RXMQbWmr5LVJcai
xRIzOEm2bt6++10EvHjU4GjHcE2t6jMY4lrwmx4/tavrWwGoglldDZVqWFqqDvcPBe92TyB52RtN
Nnx8HfEzvts/QyigWr/FYnp1788NGipKMnJrNYRZSrk8T4OrFgJLt9J8o5pDeVdUqYXPL/rmc7tR
RHVABJRqw0xXrvIF8afjQwEwNwexar2BbWWUhB+uLJSESZWqEGPphZXtlJCthLdBkb0EWxqWPbq+
A8hjdj34YlgFKQClEvZ9LKS7pRuXjm/j3xrdXqXU+hBEZTADKglsvT5wo+ve/xDW9EIxQiHoK+At
fzwgzvy/SrZJN2w8QgPYKjt44EICatMrczwbmFexXC6W9jjaaHow2hbD+8NSqi+51H1AnzSh3lfV
rXh75F8wuQwKaLjzlRxcm0pNKNIlc/btYypPizvL3kASt1T3GdeaIXBMn8u30MJ3Y2wGQR2Z4Oje
0wGfvAZddgocZYxNySEpajLWkbZCRfDAYJhlOFYRM271ekj99DSrUcPwRTSQ1LdlhzRudoU8XSj1
UefcwIv4VH4wKagvWqG0gQ8Og1B8INkzqq/Sdrdask4xsPrIHwIcjM3SZyJtJ1o4nD1X/L43ecu+
mcpTWCyuybw830S71SDQyn2ryagie7r6QMK07lhP2oK939Vd3M8vvW0yDQ0LQeBTAAxrG50SUutX
tvPnoSZkWYvblF8cZxdEmNnw/kOuie5lz8wWqsVkVs8qlzYtsX4/DakpHN5HCEfOVbKgsfTIds3S
tbJzNYh0+zYo+jSp4504GDd9AROSM3i6grGTM6QFya27DZC/wg7PAFEbrNmvzSoS7eQ9Da5qSFlE
mJnSUkWex7H+sfbHdkmbof/XDOMMiF0jRHgeO1ltb7nl3Jzfd4JEZiXPf/nJhIH3npU3rDcMpOZD
fcmz2eCDzsGFldlELA1DXgldqOckniJSgDB/KgqDlfSiOKYCC9RBbUL3jt3TJgUa3mp+C6U7+OHp
IltOj+eX+xxjOLd+790xg8YLPEOtCtR4VyG4/KrKUZtExVkkXG+Z7OpWDRUg2OgWHCuleSFmh9CU
hoHRHSOQX+MTCKz9Y5XboOsQUsJcD3ib5GYOmkazFo3iDsRb+6tUaD56dwBMr83At+rA2S5UCeL5
15kgGfa/QmQPOUuq+wkDQaCeMvS16i88D/sw7yVP/hn8RSbZpOhbbKmW903WDgZfM9Q2SSUD22m1
jTbuKaRjhdz27hoLxksOtekSm4ZdjnG6gN2KJRo2bQZlOiA2VNfcRqoWbZZ++1JHnumPkW6QD0Eq
Kxz9hjgbghFmSWWsofMS5YHY73Vm6CgRgV/8s02ugyzv+EGIwwBd+Du5CQz9fzvwppjbhGpFbR5K
tgmf2Yz4UpLALX9vo6PYwAahXudI8+ROVYo+BFQ54sVXCCCAxt2xgusqhW3iR6qTk/xQmZYpCplf
NILVbFtGb2+kH+ao+Fsr6WVAy9GK8l2NRa8/U520sgf8vaufWmj2JsxAFxtMWytBNbniK10aFERb
mQCdCNZCkeQnYfBSjZQ9Tf1F12ZlGQKOlfK8e5nIwCWbypNkFcNvv6c+4Ij/ULFfY4JxcqJj5mBh
YnJT1Sszp71N7BW53tcupBDsVN6iuPBNNHBIOsFGS7oIy9EtWtaXGYUNMuf4fUB3F2Bkx58DeQS6
L8LXleelz0rOwOnNM+Eidr1G58NKO40PXo7TqFRS6FV5YoDatFVjzSN8EuaJj3B68QClLjH4+Zkv
QNItvHBwFQt60fCfQJ6djpgluWJmBN8yjfsly6gjWv2VU19mINY0SWaN5Wa3NVZvxVZEYV6VUtZj
P42ULBbmndOsYNhn8i3LokwJ4tdfEaV1FDU/Aj4Pkzlf6wsoWktpZxCy00RaVX2VKdLCcwBOmTLg
C6ikXDIOH1FNiLTFZlOTOfn6QnUUuv0rUF6bwFEOT4ROHj0djWWbIQr5ymByJ9M2YHC1RUvM5qPL
R1XRDV9cljFjVDVQ4xTCFemvTH/2F17xZYvHOb/tSU2EceLx8WhM76xFPG/JdkrvVkVePfunxvKv
+ES+MBf8dw12KrW8zWJ49QHvIk5ECUSGgeqZZoNOWXSc9iJoKXefpqkmojI+aZTC0cTkqtUwkMTX
k14UudhEG9agh5anLlpd2yeK0AqL72ZVpQsm4qi33RjCXuvIjCnwCa9L6j+vcxjS1SMimp4KaBvY
FSZth6xMhIpAj2qOENdvDqKdc8xVRpAphwVjZeD1qL7dqXOJdex6kimc0pdoAt25c8MZ0jTff5Lp
Wb6PEnCdEE59+7plDBz45njPHjl8her43JX5SFvEFWGaVell4QfnfHJXpMLFishA0gXMqqjh5A1e
K+HF2nqnFqh4HkEk9UyiB2TUZ2KpmaDiBi2x+647DyUME+oTttpYWKpJo6MGL4uwRV51RXPhcNrp
oZHaDENw5XnfKSuH65FVBYrL0ghcgvVIErDF6/FWg2DJNPLjF0/CoFBqs+695MlY2IH2bM9DOsde
b6nLaU1MZiyj3txRMDKQbHMfZlOU5lfKboWnmOB82iuT2zncEEJVSsmv4UblkbdavZDAOgh9+Bm/
CkdDVK/G3Xc/6WIRQRLefEefj37+G09jn5dLbnSeosXKrW47sGthMTRSIpsMa/fo6xBjo+CqUtbP
o0WuU9fH7rWvzcgT8itxyDjynQ6XVFmwYTOfZgDGHOvyhap4/xdYqgiGX+2czEqsxksQULY8g624
FVrx5jsTijfIBIdLxQ/IYprrZx7M9iB6pbtgzgjuIk8JMe904IFfe9YqIyOW3SkWp7/iQ2NryA2N
bA6JBfTBuPGr2BNkx8I8E/PLe5cWpDe6dULDTh2CYtiujVZ830etPsYxuMoajtKn87POyCOZCsGG
wddXT5VBK4Bdq+MtD3aXUmILiFgHjrRNCfyMSNZjFo36+Pkbdh1QOSPi6m2/4l5pGTgLwDtNW7qx
2Q/DTX5a9nzDx1+KElLSpkPh+G6xSWcvFWt6G9R2Wz9h8uL7IZiGHx3NqKsQ1KjRYG6HmFY3hAzj
cUzVNRbVC6j3xtW02JhOIC227uUXIbiP2WDkiChKK6+alkyqdva7jrNMJYb8sd/K52UACcgaWDrK
UBh+sC30fIkGC//BTeHfkq/26Nduum01zbCS/rkf1cXKV+dcpo+PYzv5Q3Na3TephObJUgpLvA6G
XPyzUvQnpzyFSfUjQpxEMC+U4i0DmsGoBgAZLLRG6sRnkOLb/AivZ03m7ZjyNyxTiJFO9jL1hvFm
PHAOk7GlI3yA6ap9oN1F1amFyqoAE4gTpgHkOLT7eI6OnuFzm+HKXP8ddvFMlr61UbQB9+hnGPW+
luSLDSu9rfMo2rmnUV5MIo0qX+ZDBh3nLJsOmxmWoCMKLub0fXvt1HmcLy49cq/+Wh2+hGifWhTx
EXeLXXnZqFxDlsxB0FlCEVcJv+4O/vuW+ROk2MJm0qg1mLgue9S/o1fvKGsU6Wcj3xKvNHWHlRju
gTfBqKYu6JlfxeG0hLuICLUR2EH+fLV8c2r/dwEzR8oRE94wbHARuD8Z3j+952+hj1zT5b41yaxc
0c6FvGEbtRBVgGMpq59SCRChtOcACga48B0fpOcFOiNwvER+IT+A2iKyy6PJaOyOwp0rmXPxrSyr
x1ytJofFPJyazxTmi8K3ac+CY7BW5CBma60JXSrKFektZ76LTAiqPggKLxan/qCkCt8S60ZW0oft
Q6BACfLWBJMnynyt6yrgnOUsqa7FquYp6mLgUL4mT02w6VZdFu8otEtu8NniD220NNw+OAmP+piK
AvYIvNRBnE1vGfnuLB10/+b5PZiDmpokllFIWELf6Fg9vimFzk+tQtB+Sm9TnYZyuYv0JTdLRxnV
l780UXgdlW0uwxerH7rKKxgrAQqdHHqtXt16GxrVf+v+jaUNy9MsfxQKwXpS2xJLaC9HFGg6SqUx
PkigRIc6zQxg/GLMhxnB7fvHvWHPgo6JQVbhi7j69yjOHdSLnT5MHkaafOX7TaQSp6+f/yvSyxCz
qvvdkFKtiMGz8cpBw1Pa5fYu9gWuQz3plxqOjJDfuONpjua2t+HBo381ERPCX7s4AWi1oOftrwAG
EG7TuJgF78mN+eR7g2D0zhEno/qdwFGmb4P4bupUL+nlClBhUihUFgBIZjQw1ZNXg+LbD9DIhJRa
kS6q+RLWFT52OV2iPMK+9kxEAyo14mzlTdGkSpH2IiIy8yKnoDk8MSROO9I9fDd2iJ4SREmIqwlW
Nmhojd1ReON1o5dJ59+aXINSzPQ7bp23xvaY8CSutbQwfOAWUhXhm3YqyxHRP6YwzALDiYmUGzP5
OiExMDLHqe4Hbm4QobHpiYIfbLVdZ5oBYhPrUBifvKkMe8OZNr1W+/5IqkeUOxpq70sPWzzwBO+E
+Dv/WVfuvZdcbZw/WuunhrjIXxudK25dhGn56lYCMSG4ehKLYFIpHGtTk1OdANr2eLWsIX8Tgj3z
1QD6NEKUt8Qk0r+CdCzX5z+2ny6ICoBGDxgwWXuKWtacsHlkGh87KHZdt4U4h3oY3dAw2yy54ayP
Fh7T/LolZp9klgCF/OseYxOffq7QqI3ndtb75Gtryp2+n3jx1VsuS7FLLLQhbklaV/ngNS8zAEos
6SWCTDyvA7/3FAbSWyA6z2lS/1PPig4PayEiOU/Ej48ndQ7VnhQnK153a6hUbv2m3e5aF4n7BCxe
twhS33P9VX8BbmaMVBOg7OXfy0GHE7ZjoCHDImxKb2NfcbAFfhnWYjH8aW/+L41/dx6KcDawf0LR
Ppwc7voAc23vmWx42hqxUXhdXY4txS1AXhAYn+jXEKXtcJHrHDGzjGaK2ZvfkbUm6A/vtIw8qwpR
qEn+c7SVr1W4Vtn9TyxutIiVtz0LHVC+g+/lmvXnrSXal/dnk7xUhvWHh6oZjB9ij7TsnupySe4h
pIwzeM3QA69aX6U+yXi4l/T2Pn5Zj9EYg5zUR2SsSAT6XNAM6Qdoo0q4FxlRqk4fY+rovBX+hA4d
ehL5d5zAgVtcrFKe9oGNJTjKyTL17YoTGuzpMqv67jWzqtjpVYuZPF8tIK29kaS7w1ofSI+IKGzx
pI2ZNmw7Qm8dU/BWHdkcuLsXOC8EBWTD3bx3RR8fEBYtvgYlkeHmo1Ja9+MiqEGGnocDCxSspqSp
Wk3wC8tRsCDSPYhGWdqIsyHqvOVuDQ0H5kjHpIRJMAjeMDsT4OH0lVbk1buXMWKVGZMcpg3gIIz8
+fU0BRFktICS2D2pHBc3mtw85KMib2AbFY2srAUm/rRNQeGLM8IOPZHYGUHHMrHCH9eUeqO9XkJV
EfOkk1NfAOgdPXUbhbZhKPKTqcg70LlbKXcf5oZYDj6LPin3wMImEA50XSLFbNn/RGBV++K+0kYB
EWA4ukzTLYxjItXGXs4gJoF2HhxlM+sufWXPFByk3XiKUZ+1/0a933lpGVrDikAITE0VtQ42ig2w
6/CkHeqOFevvtBRR+3DLaRRCcIsRwhOQT38TDuaNkOuGi4YQE9kadpX+mgvga8k8ujqiJ78Z5UP0
ocLfwB+GhfYq1dFWNLc1w0Ur3zMsKiSJ1H+5+ybBS7naGgQMSyQpMhCC35FyZnouEIaVh4zY9ygh
+S5bddimk7qA/Bac4P0G6k6j7OOGSNcuCMcdnc1pw4MB76VqbKtF+drtpxHrdFmeONOka4OHycOR
WxRaggIpTaIJfgTab5ydoPfiFz6ew65KFVD/9YDfOIKTUofV+3HJwHCElLcz3xWE9MYqCvpsrnLt
59q+x7plD6Yt/ELlABQJa/OcizegA7AIT6BdKjgbixUsoLSy5V8zEuQwFsG67eWR+2iRtgIGzKcn
xfWLgrl4qjSioTcH2rLeLE1HzWJi+M9RGLh/kFdGrR2HlW7t0fdcLvQgUrqDtgz618xWmX06dwwL
DlVWekihJ//VUdliul18k92/aJgVFUTEAlj1iQ3hpt3/WaN0WoCpNPbr+szaHAEMnTJ7sdhw0uko
BE63fR84da5xYusykWCEkmdiLFCdLOJJU5aDae1BT0f+vcxTgEt1MUlwSPJEwtHorzLv1X7hv7ig
RnZpHwoghGjy/MCKxTlkvQ3wQZGfzdkD7X7XU8CY0C9MClhz0lK1LjxZDCRKaIS4t92zzqnPcc0s
DaFQIqzLUSijagjDVpmbt9g2LbcQwjzhVZDs76bK0dp/w1Oesb8/LWaIoRgysKk1o7cs6iE2REA6
KdzKKO2l3sagrnALwhttbolV8N4bblLYdqsJlZyjjWArhYtMTrpmwILH9gVpHrCiT6OSMdSgyNC/
ytN8RNswzoxr2GQRlp7sC6xaRvgM9diyzMy64pywCOCnXETNxtzMpotKRyZhIsRo2kO5XC2tqm4v
IqvOPTY70hTlW6a96Hsl4DbszOoANgJAt0M6kp9yapbiXDmczpGaQ0po/Kv5WllTv1a6z/KZoeCS
4iQreU3mw/ZT/nbIIVwwYWX7GeHB31rN7RI+IN832lOVy5KGYV9YFz04nSXNZe84MXP18mXtt2pm
2zVFKWYFtVZNxZSOXrL6WK39fJ8ni7f6XjvRQoVaLh9vQ0oruPR6osKenIlUDHNqfiGXKEpVb4vU
sp4AsbxLkwOgBHuuYH2tlJ1rOxBP6xPP0JpbkmhImFnE05GIRHHn7Hvsh6pNjPH6VLDpnmP35cDL
PoPxLjeqaF1mb+B0ajE5BvsSKOECfaUqgN5HL89sXNw4kWHuGO7giD5KZG0Yc1W8OnBjX89P+pz4
Kup8SUuMIuJhdOAp4AtgfYW2R83ByNAjZJA/QJIRhYwpctBAEDrsdGWuLxtDkznKJbxcI00LHZIY
CQQ+dnvXS1w6N9RyDiRDSc92C8For8OzoWDJ3inbxEuDyCENRKx+KGGh2n9CLQd8a6Ey7gQwvS2q
O7wFRAmibTHPj3ZZEiR0qBKWTmijIsxf4T7pW9Q7S/HX0aWPwXJ3+7wDHEuLyUv4/MZULidSR78G
BNDHrIYw+uOBRl9WgyGV2rW3xmLeiIPn+vkkCXCEYKQ6Mh28SQYZH8J6mtUiRfoWyWI2N35l4lcV
SOjz/sUlM87IEO35xl1NkRX7T+E2cABqnfJTcJhFXOVK1mfh42sf/5BPvFldR4aG6zgSiIeZGCfF
nwjxl/3ZbPDLEFud17N125uBIk+8zhsc3v3yiqKyL5/J3ki2eJvT1fOO0bxhqJ78UWQ4jxr9O45j
tmceynf9h5UP3Fn/0poRSSxtgH5l1TWZEo8lr7rXGbx26JJImMNyqIOVK8gYh2hOuMEDClsc4aF7
cE/RRZWM1kBKlw/vLsrMOzuvpsczS+2iXDfL+zfQ820zcChGN5Hp5EGTqqKgTIG4j+dYiPqQt9VJ
eya8i5Y+euWuiFSwb9dGv91TEwL4Gaxt3B0ef8Tiw2cjFpLPZ/1EuvOgE3xqTD/UE74fgbCOmDAo
QJRmnCIvYdIN6V2kgzs7SJWETE9h7FDROQhgzIJ1D3hxSWAumB+7PLpWxN/yivTCWWpcflhl217i
7UfAujJompDWkJ7ruhptC7y+IoEA7wIegeRPV+HUhTlGAK49IVyXIxmqBHmeOZe/5YOG0TcUL0Zo
QzW+ysJCwIXYaIn2C2oRvIPrOnkbbf1Xt521FN+uFlVnIm2B8eurToqwTKs/R0VrD6BqrO7+Zo38
7UH1mfGFFmWlwBWyY0f6eb109ug1kOEGQAL+IxN37BGf5EIE8wAWqz/7EM1t83C/2Hur4zS7RpE8
BFFXdJWIF11srP3Xvs8V41hjMa3XIQ6+4LAIRLfxms+bGsCCyE98Zm7Yb4zIo9kEICDzIl5a9Ivn
mClWoLzEIM1zkgQLjUFNhlrUa++xaE3eZhHPpwzkA0J+Js1f6HiuAAmHWzF8gaEM3dHqWmqUtrwJ
A6HSAWy9BUTCtsDSxEpGPtt2R3SlvT2u4Tn9wkAavu1RHYB9IKBVK9TKYLfRHDYdMHIaENkg/RIQ
cIkpZxQuKn8Iux6tEwsJYkoZAHAuX2xel0hxFgDNcdVf7DJTHaXQitbcwYsWERfa98zWASeJBplN
JhJXS9OsURRdon14WHzmVaLmgwHPP3jOvxRlDXSEP2KOkBUdXpOxQVtyni0SJzTqD6Za2W2Nkbjk
KPNkaJQhCG0Y5qp2H93pbuQ3e/GMRwXKoyruwF8JpnFxVnJng42PUojHI+AQaAxa5v9WjvOi5+19
bq83Vx4mb+oqKRDzDtton3Pcu9+2J+tbnH9e/pzV4t7CN9KR2YfFhb9dUFKTzQa5Ab5ZtV6eNrAk
x3yO5f+13KNp0suxSb7FSSAJQVlBb8P1AG4TgoKj/TYRpX0ToqmZDZdRjU5eex3tOISvjEbsB+Zc
DiJJdPGGBLz62Bm6cPR3An3vOmSyE5N5hWtddV/yACNvXOkDYTp1P30HhHfGz9btrX/l6jsxFDwj
mwYfK3B7o8knt3ZjjoNzNJoijNmurJBJ32nm1upBMAzKB+w8yZ4+FTwIhXXIK7LT1NZgLgr6tP5X
hGtcic75jbwN98NROo0o8f5BxVTFD/MVag2X1jHZ+v7E1dUq8lWE+yyHEfZcAUJosuaNCLeeooOb
F5952YzqyglGdpXZf33il/pFdZhEKSzwbTN4L2OqhUl3dvK+Wt7pz4HAmo+7utn4DDS2gn72jvOa
9ngL3FtPCt+8Kjbed08vaTObusVKaIAMdNga8fdoBLYCQvbJibmlx9PsAC3x3pGKZy1G5BA0vovf
CqRUtzErtycMQgXX6YN2pHGggL6bglI+WCMeSi5v1lkVCZI+ORiEQR2IediQ6+LYN+lMuwmag7l8
fS74As2CtN/LciEe8M48zTQYmuklKMmWmVcC+7J5LY6dhLEOQ+Jl4KtbWe9+IntkXGaNOw+21dwj
8ABZ5FYMYwTrWR+6WZMLROem258iRy8vEb34cg17yZPrqVVS6Qgk1S5qtuEWEJ3Wq9XQpe11NJtf
8C53WgYR5Q1bUZHehWB3u1lb+nHHPCOAvoPFkJSdxz1XTIzRuk3IyDDLFJsPoU/E+5hecuxcfzfa
rrkiOipRz5/03GeaiQR9pemqy/oj9pUOEpIF0giXpJG5iOZCi662+hCuS79IoWo76VJM8DVVoS/u
vIfhOkKqV0NMMDD71JK2jFcQ530Fp/RnAI0wY3iZxw/ci3RdFgm+s1/m7hnTMbfz8ne6MahGtifI
MWZ7RIiKRaulXdxai+zfwrsP5iL9JsIdR3g2muMtf3cRENUKeTUEYsgLkjUYwsfMvQKew1XLGcIr
279TG8xAALV3myDjGplXCaJ5BLWjCKp7efn+YLu7OrAD5PJGinYNcwZ3TNA/KYs2d+zofXKr+r6a
Mfoc+pPg52HO4rQzxrEsfv/um65oioXqINaII09QOd9BdwMwgJStSNc4oLghPTvK4aUt0Y1JnezJ
bHBAOV+ES60D+tiwVrTwtvPO3w5KxQO7FLR3GiXHH7w307hNkczckfrK/lrfL6T6VPTyBmA4jsVr
r6aHqRPJ9zmHN4b8IT/kXquG+0UG3D/1hcUU1EmleCAay1x2XBbyqvqFbf7aCXk14ISNJB/MxOEb
zmcpSPT8JDc0AlZh7jFAQlxMQCRO7KN5MQxW4c6OXhe6JgghGtov+CyDbcapuGYEhtrQkWTj+qjZ
YGdLsWQ6IKqjo1bNzN2q6R6u6dG8DvQAI5S1Bm2e8/Ap2uhPUNUE3M20CWocyLErkgVJT93ZsyZz
t0nPqx/wnKWYSDT35TX7roDSL09b1u42M0pOIlQuaXNxb/74DcVYz3rHpO7jIKP6tNO9Sh9rUv4+
/qzhwqI1shiDUaUwZLOZk3bHP8S/D7CUwVMzDcdu8JJrr28BDGC5iDTw/qNtXzkxElbHbBJRl2D0
BN0NlpxFWzIDLWHlE1ERyIG7qfDmrlQGb/24sI/Tg06stjIA5jsQP+owm8ImDdGccXriRwC4R09J
o19HuiJ2zq2nBG86/rWzmqBx+S+4uDjsNSMIetnDI2gUEE5JMqzAPe93PSNx88QDLHrlYkNvUetM
Fy+tFMSYGZPGl6mJkJMjZQRpmTKmOXSfPrBBT1TOVeva7IVovp8pJdbAKWKBUYTq8ZKzggmB1bX5
Vzcn/3Xo9gTBiJSJN9wbUgvPsxpvd1cCRP0abmv577tsFpbd6fSM3zhS9iXEzxB/Yy9xJq0FV2ZW
fUfpmyZV+JBR8nJLJ8bOEvOUAzdn4ei14fG/jrVwQqo4JH5iPRxE6ZwQURrsSpJOmllnEd/jvQMF
t4n4Qty/FFlIJG+66obrYzgq3G7TeSa6jV246wf4xkmTLLHvIRntCECoBB3kcEjtNR8veFcINwga
c9jSRqdkBCYs8KfLdAYF6ImNV4kB1DijwnTZgp76pwnYca83DIWIY+JZ6aqrIvefLJMit3CO35dC
PL0dGZEYs2MEQGmezTpxSpOl7cLBv3YDjwd9d56SzeRITs/bLx9wjeqx5jLPOca4qUuPxGJv5tAT
2iWbddh/RaM2VNhtwYyuLgzUA0vsrELw4qsQs+98Gjhy1AhHN13l/xRJZsNBGN94rjD67DmThbuD
WkM11uRzfcgUGNjYf4gZxFBlDhkmMBvc3+V0jlTyc0CXh2IjrYz6Kl/n+d7awjiKU5ocAFBhLm9g
Lbqw/Bdjk3B/W8/A0MtFfaTzjj2TItZVxn7HT8MpEhJrWoln/DSJfGp6y0gPzkYo+NeMF0y2waWl
0sAM8O27fCw4xDO2WEDR0P/x3hwE4tfu1H60Q7nNOmiXDDWPchfDX24h8PjWCIpaGhX/Uz8AMJuc
L6bISoZLNdILAT73EOJlAgL3lBRALHxmpZOd+I8Ldtfc60+QD69gR2zm8PkAIb4dYVhhdew1Zqze
+KCqrJIUZG8lA4zmEDpTzWAZA+1iaHcjI6ubwXC1erjrNrTcUlKH9C9yGiTHQz6pXeNyyTGPqsoj
zPbUKGCE185g6zUfzuqsP6Bra1CZXqFnRDNIlmr3C/PTgD9EEGjjEbB89FJVuL+FteTf8i5o2d/b
dvHSEE1n/ayeNLU2KSuAngVfJKZnjgfemp0nxq/48tzcMAooZ3UuZ3oiit5Z9ko972Ge+5RQvnOs
OUQE0rrSIbZifbBp5LRwltJnRPDTHSYxaq/HAQ1gujXJbRg9meUlAme88Azon63vhQJ2Li6iSyad
2Wcrlf2Z7a54oVyUaWt+gQGtpPpGrLtUF8JMedpT7n2CwsZcpy5vEvr9R0awnvBQw+hnWlM+Fz/Q
2drJKdwV/zTOSBXSiZO7IOKeyvEOoGi7LNXJYMLs7QHge9njzyzSzIm6WV/0lvYfmd6N1d3ZFhCH
6Uph4fkSnWI0LRGGjVVP05ZaoapEHLFTzoFeivrwpSa5wBckaBh/gKezSE4UvrvM3b5CTN/GTftU
vo2om/li9/EMp+U/Vd4AmtnB3jATbbWgTqPnw7C1gUSlKS5F0W86vN95n0d+xA98vxdreDcmZxOn
9LRFSV+vCxCmwD4uNKQ0E1oKQoxCRCK1u7l2akwmu3MJG2QhBofdMrme9yyzQvY3WwBwR/+9y2ap
ouRxn2h2n4JmquXuBZ0HW11c059Cpw0k6n+emfq0TPNxafW/xP+aMwp9ed5oJLGAYvHTl6D5go4D
8KVUbOP4XLnUJVBRjPxWuiUpdtyX5SrnwHWV7uefcOpHRjeNsIRHbbPjbV883oASCVBgQS3PtUPn
CbkWqHkYXf58CSX7bsjLdn08hko3r/2mM8Om36+aUoxn4vosJtC3Jk1whKqNLjzvK/geau6nIr59
7rX8vXMLuwq9oQgpVW4g+rXOP0CJYsYum91xsOuCMnsog5kcjVF18E/WMr7faicTmcbcyQQBtBKI
KQGRLcruWAjTMLC86QOrVexzwTTBpf6tM25kfX8cux+d09+4ect2fbABrDIHvsxTYOUMLrpk2NQo
EPbOmrKUFvNOf2dYv6/D9+uO4nlb2bHJo4YgRzMqVC3ZIJTiCl4JkUXrS92kdkwXa1+42HXSlkQM
2eTpaBoXPwBXtFn3XttKcUZ1RNj3NcumL4wdXyb+wiBZ46/LhUIC1suoghPDJlFnSG/0yaNZhWhr
zG+ImTEnzFTb7w7XUC7ChiVq+TXP+Gf+O6Y8VeklpIJSVgQ0fLup1oefMB8UwEAGYRvp6B8pdU7Y
dQ64taM3kYg0wGlgJ5ifuKgQBGy4PtPE83R3vLgTFoyvE4YhpGL1ZhYkjNU4q7XLGWeB8j+y3EM6
/Auw/nps699ZDpCFNHXJqXQmOdRAMRevWDIyNkAi08JFWwqSNN8SgMFCYOzP5YDocC+u2b3AMy12
/Q3WpwucvS+EKtD9JiNV5x6eFHpZzXIGraj5qxlxqP3sSCe3EnCRUvrQJstioEhSn9qPK3fcayE8
3ncyC6aG63oT1lcRWSKGouu7SDeVap4W2frg+SPV0/a/Ji81q/jDFvdUAa/5L5W8CDN083S5L8LT
6dtIrUPxr0eV/yKv8Ngwu+bskp0f9QY78orVDGk49iXDhORbxoJbqQbVxeuxZrGh2mGidfrfKaqk
YVnyPHv/+kVbZ+ojP5Ow8RsPd2tgJaD+pwKsARAMP1ltEWwdKBrAFP3RXo03gzrDXHjnpTfT8wee
kGPMtgj1XgFyOWa13xeuFQZj9GwAXMvx+lQsjFAlQaRY9NcWHr+roFRq/CmLhizAccqZmt0LWEhO
THihvUi3wB9M3zUbuZ+4W9TEL1bDdzqolHp4z/OBl2Q4yp1zbsBUIXNpqfbYgXZS0W+hWhj8GjuS
pNr3E+tQVNh+uAcI6jhJ+b6mEO2GiaW2VOfEOl7LPZ95+0Amhl/HDhglTrYUT93XvjsS0nL5/c4l
KlPnDVzWseNOISJqDqejZbJsqYvvsao2lttJ9i+EhV1x+rooPmFNxImOSmBRdRr6X7bWQtAczdPC
Nag+ch9xyEPw1/knJooefP0JyB9/7KIJlHprtpJQb/b/HMj0019ue+8fJyI6WIy48u1QlOIQqnIO
VqFkheiG9XEpWEI/MvLAA599NmMr19TOsC9vw1Y4kq925513icNOjGVUVe+RFR8P91tirMmLW7Sw
fq/4y5p6LpI6AlWClpOc3V745S4dKRgPTDh+g4C93L0qSNejFHxJP2mTCkXeQLVdfJ0WdX52sSxi
zJGVeKEAR31rhXvIKo5Hyv2xjsNNUuFpJHg2Usu9SS0nOLUaoaPXZv+KU0jmjdG0raWeVWFrChyj
VY7a2g9nQVILGJmMVLSICTL1122BfBbTiLX7IH8fnl4liupMEb1GXHf3ns5yZxhwrEA8IUhVy1bG
Y2KbMI220RWUdp8FS0MoP09dKDD6vTIKhhxEmiNswPRf+ZhCyihd+zJVrqdYYxeJgpLQQRbAp7kf
RQENdadisE8u5j9eSUsgmu1PlXWGulzotEqg55f4/+CJBv5QG12RHWdAMhgTRiksIjPE4oFbdCqc
lsGG5kn5E7/20A06tp5p5zSjnfaV+XguPUlR+07jHVOvEzyeU8Z3Xw6ko6cWuQOjQzqYJO/bXTFm
+1FdPvV1j+2NiViHbdDynH2xN8BSx0CR4vpdmQNg2ooRvB6pHI9XI0w5FnusEcqEpD+kFc7XwTZB
Mmawl1BSx3feD5xU8Suc58XJK93jkpxdUZg/Zl6pN4RTqiA5JXzGr6I4Nx3E7aUFE1NBKBKAgk45
r68Oa8g/JN0TsV1CGE+9wTrWX4hgpYvH/6qSLL2154TvtX2JXNzxZS3IHB/YvFDrtE5H95QRH7pK
Ix3t49+B5qGF7zI4x6xO59f6nJW3+kc70CCL1Ift+mBvQHUx/tO0qg3G13eK4rJ+48JUyTqNQfi2
AJH1vsUDBkhNIRANly1unTWYtoFVS5j5y3DLX/4ptf08v01UGhdDbK9fS0dWEluzvXUYfzn6X7ml
6mnKGJhUsLwJ16h1RPKKh6A12haLjIWnbAZ/lEYEQNkXVewR3Hf0HT2qzEml62gKwZy8Suf6GHMi
6BBOk+FTJJK+sNaqRxeoi1EUnS+Ixs1ziKu5hYma688VNrh4D6B3LOUKcIfejs6P+f9tOxnhxt2U
qD2oVvQTsDkbTJasDjEJvpVh4XEYqHXOq+eCnQVWtKML9f4WqZ9HMWmttQrIdcbhQDXEGQzesEXT
f+YZIQIeRJuxhqLq89hqBneAslgBEIT/mZfZvA4Sl8qixkmFXOf9VleaKXSby3/c1olpOg0a5gbS
PtvXRmDBKh19WWZQuKahKyWes55Y3aXpX//VePD3cTRikNQfxxQNPxYYsDXtroYM3ip6hfZQ7CMN
q1MmvmdFEUBf4QocSxf4xeOKVO4UEN9TB2aN/D9e5dMgIQvZ4FFcVcpKjIqnhbmssEEUITQQUBEF
KbbfEW98MWxhI/INK+zcWOKr2duj/kM8vj/qY/8WUJ93XtIGrir/5qDROReA2cv6a8L3ZOQ4fc3K
izd5ihYeAQUcGRYXSIDuHpUpxbJYjzHhZ1j61eeD2FBW3kTjNBDK8jBkLR3mdC/qGe0Z5x+gOIzP
GNI0Rh5C68PxjYLgEwHw7kphsupwEBQZunPMjZZ+67uWRGgVy3iEbWm0sQ4pICKtxO6EXo9IqVqI
+L/z2hqFEnTlc7794vyPwHRuX8aII376Mch7T3Q0pO1aIRik3jAFnB8cSNcRI2mxL3K9EJjl6izm
KfpDMgLB8IDBtr29WPFnCGQchL7LaXTemE77fwW2M/Ul0i+zAk4i1CtF3J522+GT0VUR7vw6qYak
hjKNBLZIqgr3K2r/rYhI6OGXcDRwNjn5Tt31jlI6utRFgwM7vy/SojqtUKs8i6KO0PG7Nf3NlP1K
05kbTNl/HCTaQJmRSxF2F4BAqKUMubzqyS5aL5YGK8giN/LjZgEuYpQgLTMWpVFLbWU0SZM5v7Aj
HISa47UKSyu2sbJR6+JwjqzWle4sPBCpPa2Ek2g6TrH2U+x8X3blOWQpVpRUAa9BlcT5iu3h8uvy
zgCZ25muKLinui9ZdFEJqVDKiMpITH00cjStBRkfJbScOUoMwiDYR+DIZ21OBcEb9q2kBBfP/As1
ZIV5VzyNwb1j+VAVw+Z5W4NlalFWIhU4oEWbFEbTjWEaKOTEjiyLx3ZErsNMQ2tvqGsEmz7bvxTI
PqxpoBStuh/TFqhsOT09ivcwLKKt2hNmW6v9Abghq7GsiP8Aoeu94tmCfz6w8gtRj0BPtblLzT4A
mhm0ACczpunzfWOV9039xvcSQtuC/jYSYMev2QD2H8Cd/Y4JnG9POYtKzbgZTwGyip0uHSzGLpIN
2CulFdlJdcpt1OvNWsoFZsRuW17g5fWNxgtxmqCi8lLndBD6XMfsVovaiaFEXS9xhrvFQSleCMI/
PmHubaA5qmJ7P4pUTTnIzzTS71jOdhXwjutk+3DQVBw5qALXwo80Ol6Y7QBHgVI7ieTUow6gQsE0
s1LqSEDA92ytptu/DGqfpjSC+qt6MVAZuXxukS0VaMCd/30OL6XtBGN0vkzLm8rje+oKU33r/qFE
lp3gECTZNjbLBXs2f0CcF3gu96nRpqcipDj+TPTa+FSVKzuC/UuE+71/edXVu252QzuwtOIbsz7O
HsJtW0rSN3RH6dP/ziAJRxR8Ur/X+J+YtCVt0XdIOGXhsKXgXduacurT2cbq9j+jcr3k0dPkXR/R
lIQU8lquXPoYoPhj0LCrvaYskPQzfYMwzjvCVivo1vBTbzz05oywRD2o02Zn1W90qhXeeWGjN20K
iz0oTI9Tl/Djy7PwoHWfQCii0FcbL002mz4qVwV9p8pmmA1mGVZGIUQEbccisRLwPer+XnBnkBip
1xPDsecb/7xTT0WgCxRWHDbMk2F+lnQQG6IyBxrponClzxnhyCZnXznspv+aatCXflFNWhK99SEx
mkUc4rg1B3lV+VtvydkMihbGQk+RjQybhHQoeycR3cBom8glUr8jadwW2Hp6d5wRFjXYz2OZgau1
jIzlkOe+I9XwNBk6KPf4LSp7HbP6RQxJeSC+E8f/BjhvGaBRuHVf6njRFs7EcCk5ISUUwS5ipFYT
MQsOUbitjIdT59V6FQ6qEySyYH5UHhhNxVPAgwcEF/ImRZ/joZcLkododeXx+UEhjUOHXetLc/p+
EBiiFbJSybt/CQUXffiLP4l5RbuwO/lbcOaInXlLCB2aWKfxL1g/HAW5QKsXVv8et4NMUvLeCVTf
NmEoLJFErmiA/GmCv0kzWGbLumfLFA/StAUIH0virDZXIYvuWnk4NPtFl4vcB+x3hF7KDXj2PBQy
lnHeK+Y0xbkU1qqBnZgv7M348nI7AQZpmNtI9L5BUj690FgzoMC5qmaNOjAZDuYNwzjZeMI3z6em
qL4GMRE8y+J5dKSsE51BWE1jO3NiyMozH34viL3bPT9TpYDZc/rsSfV3lnsaNXMFdewVBIGdciim
K7Hfngx2Wl5m/41i/osFMBy8KnUwDte2NFq6U+xhJ6Bd0Q2OKvgD4jMDJulOLYirQYi2UJQDoC3v
5Ima5+l1p1N2rpDI69B+bXgD/7asAPv+VsCNhWR1HtnoqNUaDwKAWEr6HVYWw5niRuOidVong9Tk
jY4sX+TBdlPhWOQp6L9e/V0rgRYjjVagaTqfvgkjXx4gkTce064kufk5QAvu2K6UuZR+G2t5K4Gd
++wNSDTIDUkTGXkt8ZN0BNu445LlqIA0IqYP4WJwtxE8lGaYwMFYkcc0zgb15i5DEXIgkiloswAg
5Ro4wpTjx+k40yV9poXwjP90vvAFe3RqtPmJC8J48MB7evn2mkrDq2UGMO69qinT1aMn/wdyz1AA
OmeM1zi3YZVKgBTjUSCEdDv1VbnKWnycB2zGor6aEFOsG00hH9jjGRGZLIrEbsvYmoB4IhZeh33B
5lPBKDv1yJUAnKiaSMfbqhgtC9Lon/4i01lPcfwSFQ4DFCqrBQnbPT2cEIFCRcCLvbYibggDk2kT
fzVMF1O3sIJuszfe2VEiFY9itJ2SkWEGUTE3hZZbGdY9O8t9fpEy81lkFTl0YqE+l8jvZh7WjfpE
FSLK1BAsqRTox6BWuoweSpLlgD6H6RobidPHC1iZ1LIDC8df9STr0pqoCaVIEIukwxwnGYxct2dR
JMe+BmaIlnKWbINiJUCOXtQXk4cVyTcGquBEuCeiDyvr7baffOUL7GQiHOUzqUW93BSCRopc/5Wj
nphbmI1c3NJbP8tNSdbgSLOlb6ZqRyMjMdzYgEbIGtcdtFgCgHx7G0jAhYGPpNO8wa47bwAW98EY
eAKhBxy0TClDxA697GqGMs3Ce3e/is4Du1tyKda6mTMguRRGhGYtUMtcf6ozCQivoVR1UFboqpNW
WBqrrxzBpgOfqE7A2sZwurvZwEvBZVfPLsmnHMBWyOz2I229IEpLcSxsm48yEMmsgwXAG7Ogw2G3
lTlcyketj0wWerBmZaHckAGt3lXt2T/NJu2ZsvdpESgOEexy/WgzmjTtRnQKsQZGPBaMSS/yih08
Lak7DvbtbrD7hH06NNLBKIp9M4hExnr29oAc75qlayz2+OTdBmvuQdU5UzoBj8penkJDMXHcnqK3
Xdd3ZrcSM7UwOtzgomHoE/QUGxpyvMUbsZxIA/5KG9OcmWo6Z8JDS8fzTLm+4uzI/ldaX0lFh7Lm
A6f+WsWwTXkqokXhxKBvYQH0+dV3Dv1aOIXzDpYr4CHFdMgj4nefQXTRP626x+nY+97qG8sgfYo3
ByVHdRkcvSX4/JegCE/JbSt5lxLaKx4aV9aWF/vcnpDsFt0mupk9dtKOrvFhGXMDkq3LGzlGaLnE
2Eb8IiCQoBZkdmCyiwxP84jXbQN0sJwyuTzt7J40IFz3WRixZB8uSPH2vmgVUmSJ323XIvYIPC00
WP3p18aG5uaqhmJ+vsrv3MxDEYplp1y5yx03OBzxuHBOz67HC367JHO3P0/mNpwmdnucoyMfZQ7z
aI9/PPFx2Km31YsQknY0B19r+qOKMcoen2qPeteystBxkIOsIwAsIswS5Jw9AVrjZUPwdlgI4cTe
/rdCkCmkoc+9FyI1P7ffBcSTcc/6CIWdRFPiS9W7e/nGLfvl9hnkcn1GsPTr0gh0ZJEAqfURZ5rF
vgHKRYCRN803e+LCNVzYcRKNdDUbCIcuA7VxoFVT6rEDkuXlx/WYwaUbF2NexheJMBpkAEA1VlHP
obOnnF+SwSclpfwS9mG4ivTuTu2B3rSDkix4m3LFmk+8FAxx8zDW3HXO4FdTEzLK/NXiHcGaC6jT
WzANRZGLfUNOrXn0xRkW0TmyZSa7vkeZ18VbT4wXz/UJm4ZtD2toBbRa5N/rWPRQAbnbBY7xMY0j
h1GJf8G8I+LIfv6v1GOBiDIqlIEEjDswp/VYDPY+Yu8IPLQOEFrBW19fASDb78LqUAK5bCZqCSLi
fjDtCFofOb1hsXcGTMhpLaJlThhmLe3H1ITqEWqSRW3lVVr8ZQPEseBcgVe1DI9fVukcek1e6YAo
TmjS7RIDD0v9V5TmCUAGsSJSbKaQlcuvedQK4V6PB00TC/jmk15AeoE5zpF5BsJJ/7o/Cl3WHwQP
byz8aNhZ5Xio3l30TycUrY7zxw6Nl70fQKANkt+kvgJhUs2roTLVVl8NUry7TX6XGNrs3TlPvmd+
Vx9S1gtU7Pe/5UEud0PBpKfPH1Cm+M2KZwWBIfrGDBVGRNVbDtb9TjRD2BgIq6Uceamw2PFNPKnn
QULeOFeLMBeKVTB0fkuHiXauaMcvB8UG1OYqs1qicxSqX0Nggj9FaXiz5f8H+xgA8vmUZMY4G8uo
FP652RahHTbyUhZZ/yrVHbyG1hmZbfbcZ+I4t80tq+OvgCU0GIUaywq38KvhkRxyavyUTR6QPRHT
ugAZe1QZo0e4VwrCZwS1MyWNQiAVCOAsNlMrdKIJQC1f8EmW013LHhx5R6gkwMryI3M1zRNm6xVy
tSoSt0gtBSs+7jTMKAFqpLkbWbUfRkrN+QD9OFewUp30PgSWgeWRMgqsA2xg/AXAoPMqVB2hsmrP
K2muVmQGmTzfNVDP4IwA78Wgkezu1mT0utxW0OsGZQWExx9T8Ov1DneM5eZhM4yhnthNIogXjGsc
zwlYjXmys4nWOjVXIfuiw+BiJsUq+/Qm/WW+lLxdDNT9sP0iUum4mO1E+OhIvAc1ggMZEtiCmFXp
lL1U9L4r/Qx1rbxRuh28XasQSMCUTIl7GcPX6EnEt5FGMbaQlBL1wn54GUsnC/XgvKH3IIP7h63t
JLMa/JV7yBYzG+7ovGh95SO+dmbdy9JxqVqbzOamqqUjheNpRUFkWbG/5tAR+35a7MRmfogHbPRn
lK3lE2A1v3T5h+m3ztmLRUeq3PGOVznmPpTiIVkEUPVHsmuBSf9Tu7AbeOp71XwHP7ORbP/qFvXz
3LvMLzAeXdBYCqp8PS0qYdBeoAIqKtMXkscg6SUy5C/QHq98J9stZCKVe1nV8jUhrfkCBtFYugEa
pCS8XLhQ4+Vmmo5De15vcuRA9eLTgTT+1TqStxQ7TNuNQNvlzJX/zmKkywafIIC5veg9VaWIiYwP
euaSmcHKg5njqi54f5g0ifc3T6TsD3p48mGrVi8r25sEI49ggNH9afdohQF6/ctHAqh8+Gt8t2WX
meYQen2dCKRpUM1cr3Ouv2RtCDRqb49ID//hE+DNjNmpvClIzLtkCd1NNIxX0iqwajcRbqEmKi9J
EfSUuTEePe+cAkW5+Ad3Zfq117MUeGbj34QBPJE1CM6rTRhOFGkD/oo3bxE8pkz1CA47VUZYGHme
m2SPFP/MAO5oyQyf9hczS+slpZZcMdngF+XHo4Zfz1Gp0uobgLxI7OyPdNhQ5qZMxl63Yaa3rz2g
9sPCfsYOxMAz8gQWvjJ0ms1Evi4YJd0L/rJW0/ra9a0MuoBPYEBvMHdHtgnsCLyu423K9tQDV/vC
wHPXPaEUCuVlxyQTyj/YPtGKCxUtLMhJEiZstLhRhhtcKQgr/+DBU0TxJCCiGp9NpxH5aJ0xsAKc
Hwwc8RJL7dMJiu+dNIgbPFjBO0vaC0uOX0pmn4SifQI/7YoP5Q76ZHnXTUolmOlbveR6d2JlwbFA
fhY/tT0vAyuNsvB50M2ArwvbauUAmn8FcmFqi0Rz6NWpx6A20b7eBofrlUR0FxllsSDpb/jG7uhr
DNyIR8OACO80sdUbNALNjEkkBG9BnZjGVchoDGLLWsEkORQR6veIG+QviEoSWZDty2ZqsWvsHwQL
GAxBQCUDZqnVOjseddxbvaLbgrCfNRjgiYR0rLq3hwZKUQpKXj3NoqVrt0VcmuiHmZlrxh4Ig4gy
s+5x107DPjT6im1Nt2IXDP9bXTB1P7e8HEn0LWSWXxXKdpyXiKSlN8KHmoXHucXhHK0QS1+PRXF/
B3TEzmodX63ZwHFXNZU3jzSeMRS3KXZVJ7XqX+tG1SW6lRHOnYWJ+57Ky6iwZwmNIWLa/WZtxih6
LTrMkADkgrzNzI9LXKcIP7ZD870e2EmSCMOxcXv4b+DUB4Lj+WRb4R3QvlUNkV67ixhI/0Qnzh42
vLiGWTbT1f/57BUrCNZppGawVGDMdJc/yLUQKVc3Mqmn/t29rY6fOuWL33RVBx5GNqE1u4bk7rqp
rA0lNRu2Kd2y3S7YpHH3n5yBK5u5fPUXDzdYckGgDBuxjegMonhdmqIgnPz2wnIBUHp3UrC6CaZv
JLN/6YzOLW+Igsu5c+YNEWRTRapKkom7nbueNQbyPcYLoAlnX25YDKmw36QDdqEIlrQD90ptFvkE
RE7xTSnXuop7ENvvD1PA5c+HEsqhogO2U+ZV/Ahux3DI28aTT7uyQODixWApuQ1GB9V2S0L9JxtF
KumbXvQ=
`protect end_protected
