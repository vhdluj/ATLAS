`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H0ygP4yS7RPIA4Xj+m4gBtCyQgIp4cZdSLl9P19Lhniw7ZqNIPGSmnvWJQ75tyxGs08lBNstknu1
ZGNB7QKmHA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IvGHLGVpLJDDlatDIc7qbBdeylVdkaoNyRXJvwXSjD/kCHYB0MmwOtDVOlcD8UHgJ5EK9dSSmQvk
H/3lSiEdJzyGT/GEFDCFl3zb2EH3d4VUguY2JTi0zfO2Je+gry9H3MgnCXkL3RNew/4rbVDG5zce
HHFlfKyFwtzjNOClDM8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nBCxZ9c3McIBJXrU1EUQ9a2Ngl8xz09sT9TE09e5IFNsB9eWAGlbChQi9IjHeQ9DvFT8jKuXNxbF
cVgUMvfv02uUBmcxYQr2BOb5XcnpdThQZ89+OxhV27EcefnBOyR+OjJm8NNH0254itLIY6/Vi23J
QFlY4qUOJF35vSyl5W0plqBc0Pf3Scq6GAsWXiieN765COEPLEismwbdqoSgHPlSfevxFNiUwWo4
OxIVeq6ALkGQ7bta5XUqs9Mz7UnROzCNOFKfRtm/eUgUKEErSQCbi8Fys9Ydcdp2BzHUS2y9mBP4
Vxr7/zGJp0FKsRQRkQOzYyWYF68WY4Xc5fQp2A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PO+DBo9piHyGwMJ1fPKGlI7FqWWvRn0oo9vnbmncuCxMrBEblZSciZSYObAah2gKIisig0uje7lu
tOSo5hNuyZrsU86hRiJG1BsxIi3VbMpzYX96CMGuCotnDOGdXSWcZhot40BTjnlA0dR83Lb3KlLx
b1yN4H48oBARFTrlwGg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SYM0yM/z591E2Z3PR5qengvyEhsENHJ6B8aV6KJPniropCzjra0otIzPddrvH/eDJWUPLjnYnUTF
wl6lA0Jh4knxsf+0Qx9cEs+wyhbVT2c0gq9r2XrjP0RJe1Az5W7WA0tEfMVv/Tc7NbdpbnweZKJX
+4MnIEJJroZ/YpDLksctXSj2g7ThneMeSoX4fZQuqtxUqeY1zv7tJDjU0kwwdKCdvq98BmriTQZx
TpDf2PErHTVFA82xFDmrv8jQqgyK7TzzRgAPpWOH1lI/gQOWf5Z4bpaxs2cw8q7vBxjwrZDiaMsw
D/qLxyw8kM0GylRGMbIUjvBcDi5EXFBjVq7hig==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 27904)
`protect data_block
q6IE0Q7J418aTQCwiGV7lRGx/Kbo/cb0qsgnRtyQTi7s5ZRy9JpiImLa5qUB7iYNxulLidNLmtCp
Gr+Y+LBGkfn/x+Dqz4AKDobSMJhHsj9jSuySkktEhD2ySq0OYc+JPnb1w5KvvIRSUrjhrbuQcEOm
Ux2Qdx9PNHbz0IP4Sb+sBtv+fZ6VwRvaNkTgu+KFkhIU/kaE/uvpZNP02vJxB5NHEnDmn+QYE4GW
YzODJjQuHF1X5xs33BlaIE18UvgV+hszQ6VQbJUH+22058/TieF9MKoHx8eyoCyJspY4COGEQ2/K
h8LCwLZ8FPnZXTgrjlTBxISytf9OoHbe0ka/yTNKl04NoRRDtWO0vlUMsHcBptxONyimmsqJ8uK+
z3fxXpBIk4Vk9Wn7Oz8d8GDcnnPtrkNH75pm4HLuqGxKbIs+c89JcHSWgyuLdgbyx41A2/bBGyHo
Ca8jHviBoZwpcO2nvwSjQ277ZTaBRECLcpSK7RJmKQdpX1+0+z8HUQ3ckOc3zxDXMQI/rSyIxKQH
yw+z3ozqunX8uLlNrQqQa/9GCMl4RSXx9Di6umlsyhpjLlNv5jdHuRqOQ/NyKBTBuTIjOGpKTY/i
NIHHKlhDPGt0tsRTYCzywkdP6c6lQkjpAZbJVjvfDStCoTO6YQPCoOl/05pRGZYO99xhhQ1KbfrZ
mwyy8oPaA1j1rM3JzxitEKWnRnnVjcfOA++UNg4AR0Duc9xtF9JFRPYwe1jaAag6EVrq9L+rb1hh
frxFGVHiCx9WyUChfohlMt8xQ8EykJywa3hHjxNAyzqtGrhGLRF6pmtD3Q1lovBn4B486gd8Eref
o3X+PcSisfofL4IJJAYnWfpit6sqp6Tx8keAo6OyAAoPdOk0dGlTM3gojszy99aJpM85m1ZtsnNY
YaxIe2XL5fNKJB0wbDR6pLCfV70DTQk3z3J2FpXAvnk+dr9NYATo/dhlRfrJ3JG7EAD2iG+3z+UJ
MY8jQldl9KpqtRGLAjZFHjvmTIO3MaQsbOUxXd7sWrxW56ZxHtN1QlEog48BO6chksniOY068xLH
C8QKUo95IONKMyhEi3T3Paenf1va0N3RmYYRihdoCoQLB0rYQ27PSmQLZE5ZLkMeOPfrKR2M7If9
qZbNjI5Qg1L8C7orsmICzId9fpWoNxKTQ204M2WFhftRJBFz7MnVS338kcr6zp0sFj4Cf54oSwae
oQx40Y5umk8X+Ha1geegy3TSoPq2v04NkI5u7fE/E2yiyDd4fKHpVyimQMD/r2guz0w7HherVlBb
Zta1nDJGUfelaIo/0tbsSiEOdB6ZEx++VYmeUcoVlaCywhhwriZINDqhY15bvc+2DINpCmXGEawJ
h+1tFB/+ff7pjT+RKTkEbzkC0b1AbjBr5g1+oJPwtxVlONDHo985TCRbsXd4P4rhBKSl0s9zu4YN
/+vgunmLSmN17pksE4Qedv0LGkdb+k4V3sNwPaqYi2RbkWtOF7XGzEVjGqr37h8Dy3cTzw+GOn+L
DkPTfd0a5nSuFMW/wkkKRNZcqU0Za65X6gRD/wpoEA5nznx69lH7WGs1UhyWPatPurTZ7eLi7rj5
Bjy8a4HdbTpr+EgQqQGZI9WzQ9We75S0DnjUgKhCI0LOdEKMh5UeqwUM4PZaPgoaQzuIQGbPPoQf
bRftFAZC4O/QF/YNaN2SEZzii+rD8gETOCxpLLckX1Wtc4Ofv4+lOCqRxIcvV8205w2BOjFnjqeV
wZlf2MksLOS1ZAaAsoUp6AHlWnyGsQ2upkP6Q4A1XiKpwM6pQH+Gv8lzcZgku3chXgl1CfF255dN
3OjvIYCicUh+7tgfbALirt9VRFObZkGM+hKIiY7Jor5lvBp1J5Xwhv6wDtVRIrMHPqyI54FK+DEF
PFRFEk8YVtBLtlkBAT3w0FgVfPTgVCqgm5vjn5T37AqPuyraBftBgvF+wGccjDEdWu9Tul4YoMoo
gTMGsJEAyaqgBJN/zAVjbqr115J6Uza02mtk19w8JPiAXGStK2i4mp4ejuJ/zx3RCckE5Wns8RKd
00SpGBZ8XSxpkVL7Y1u6pU7g5VG69x89RiPsdSEQZFHQm9mMFajeJuURdoJcetRnKt+tWpvqoJo+
aSOY3DnxO8n5xMTuR/bOgHItNfAZrM8r5O+cTHM30Yh1KB3GkeL2nexT+ycFI1XHJAtgGr+VRgRb
MC7YDQP03P+aKCEfolFSG+N2EaZDT6LTWB/c2dKMEsMheNZqnqZiVjUeXZPWmQcsqIIrwakbMkm0
lkapXPZPId0vsntv3LrpZqtZVe6a+Gkb+2zSRC/VfaL424bbF88IK409cXp10m97PSwvfFy3oYYA
CvxooQ1bZ2oZkxz8WbL/slNx+aQWcDGJ/pn8HpeaUUQzTKTxm0fNKrJdG5kVNMsCQGZHkQ5R6Z+k
OiQeIwbfB1DmeWXcbYJyB7rPUkinPIaAjxvcy/kw4/4Qu+s7nW/lLXp0jiu+8IJsuNq4rojCBiBk
f7lhXCk3zQHLa9m9Zf2NDvHTNv0kPsYH29eDF9Ltu4GdlOH78Tx20yICkCjNafQdU++FgYUVyhxg
vMyLWKyNa9hnvM2yWSfmEB9pburwXesNm9Ss/YNFfZtiQl6UQE90unzmnrQpH0MrazShv6FKLFuf
+UwLMSSvt+MNNmUDncZPjM5TUexZR/eaFvl1p90ThmR6VaGl4VUsFXeSm5LS8qS0NcrYhy9a4IdC
IKMfiN+kMZTVstJ7XhUXz9/MF8wxT1ZkuhC3q2yitOK1V1nUlvfAmNZOWfrd/j0UDwbH5JSNSTYc
kkxypb5Lcw+p9bnIG/qdqElhYVApzTvfh41nobYIRzqjPnbVXARCdZW6L8Go+2Kqshw/VoJa2Orf
RhLoFrt4daPTs3Bm3vndp/56j/13rQTBb8kDycJkU8lgW/KgCyKQCQaPkhZvT7cU5qAOkXPSaI/G
gZ8Jq0QInCKE2KXx4XifAonN5LrOBaKmEE83wyW9l1jnugzAWziJla0IypnVa4Ac+zH/+Xx+Z+c2
EExeoFWWi37mQS8Vp3AfJ7yBsqIdVyqUmCjjOR5rphGOneZyfxAvSSuKlAMPuGKsBnTCh8fcFXkc
r198qMZbMW5ENuAE2SDjlvf9aZozAHveYJCm8dyeSGt7UWIZQgMlu54bniODCySArAXXgVrZFFQs
w/v1u4jR7rXX8UyeOlhAZpi1O4bNdsERj9zQV/Q15a16ACDRZmDo6yiCTmepUJSPkiJ7N55xb9Sz
DvhzruWPjIhWQSXorc1t/CW0ysKn+w+bm5Lvboowlj1ICqyKDmUbgdFjT3j71SSjJ1+waiPkT3xY
MN6IN7iOfRYxBggL7G0D+kLabfU2B0ENPLiIDK951R5knZkp6FYlQapYt8trrLUiEip5v/NPU6kY
BmyG368c2IUy6tjk+tKcIeHve3HkR8e3BG41DfLI57eJGh6jE23H7Y7S2kFq+R5/RLmx5YKxGDgO
ipmn5Zx4MHT9CNsEsL18KuyQ+dpxPS2FCcLImRnaM9SH71SXcE729tHO5rKlYw3CdtGAn6u3N5vA
keIeK/YxGP1pKSxZxlrmd0oLUlPIxdULtItvy66hcGSdWwLw7HiCGp5UksW1tsG7h2RaMMxN6OuV
wNo4qMGn2KuXKLIN0fWxLzaqLWbNCA3Q8PLnpEwLWxaPO5HeMvRMQvl2k41kT8zxfRnfK1cPPDjS
hf75s8s3IHwWJcw7jfUFRO7ynFh2ZktaOFADYQDNzx9WG/X3UxQk9DXurUO18u3vZ1Dv0OmRSpVT
nwF2WIKa6gqNqjK3PTAmLtrRXolKX1DilyQ7EWpqmJVRZJqSY5y7uryCXf2jQNuMp9hF8iiRVhlI
m9/r8woOIwC2zgG1YE11YCEQD0nEHwAouZIUaUw7uTqnBmcpqI1SRlE9rhS9xjZV8UwPIA0hjC+K
7wfyKNjK4rB9lI8v11Hs9DEtR9zscSqe/MXBy17oZAymfNiU7IfF6ZhAXVQelOyHLTNRf+ospJtP
dZL4f2vCygz6HavndLJUeogDk2cr7vzcH4zRf/4xDTnLeRF6uHV1KOw3bZqgQO1YYzbakLuN7key
IdrPKBc1O+eKVfl0GuC2yAV4pY5iJvfGEhSpmtP+RtfaYhQWncb7gNTThzYAU05X/ts00VnV2o8+
mwYbBTL54kRLfCszKhu2XsvYK3lHUuQaYuGlnKHxyaXS1PtySJDhNKJL6o3VhWySURdc6nylMxWH
JLjnRNfBJLX32KkWilHAYblgJ8dkdnXZ8xWPVYPpWruC53YZDNHmhV4jI6NvTJtra2UGV+OIMOX+
VAnqDe2rGMnz6bkJbcqcSOyE9QC8Hn0EgqcLhr0txw1xg/UyQNMIU9e2tlyzWl/Q1rxF6/kqk83E
Trkr7drQcYNGJ4fSkUQQg30nekmvE+ECmvIanag7CR79BG4V90n7rnnR6QuxAFF9afeAhsCc0W4n
RRqLaFaymBVeKLSguBYypGM/XG4Z3JCdhSRTg6LaGywErQOKvmiww5fQQRCBJztR3Ib5TWUz1W6k
5uVN7hn7E/bZd+FE2wA46WvrgVFfy3g0vxN4d5psYwpeW4PU/l4uG++LsQtOkA/CBeloJMpgI8hV
zWFLKgeSr4FyQYRPQO9wmKthPE1rSoeoS7GMt8kLfWgVi66sQcheDV6fGvlZUIYB6ZO9yeXAxe/b
2ZeuVzcKD+Drg4aWj+k8AM3EprSKKafoUziMkQlEeXefpmVwkrqzZQzVabbo/RVv3VVyClnt7TPE
9l8fQAtAVDPY1AG3lS8zvhPGVz360ylQCsrJPUF5pGIoYFi4hfpLQrDnb95zMSYVZ9Z5qhSXHhJg
jGkPU/icV+QnLo9ih5D5thJEeJlnydr0+ZYqxcSiz5cajKgPdi84ytfr7tn4NdYOa+7taErNNHP+
yEjuikIn2tRRoK+bmjMBTnZYgY9CJncOQ17DCaOQlwNRM7JPVioxl110QJm5Y8KGGVFiN5iXcLYR
1fA/pXWkdWIVjmnMNpiuMS9Bk1q3SsNUjypNULMTpRudBAbz3x9Hc9xSO/9P/TJMr5fqkbtbAkvy
n3uItbdFygap+m+74Rqg/g8+ycwFvVnCfgaLaWZl1eYn9qRUlDeJ5J67+VHQ5QN4Qd44F94MbNfK
iP7r36XaLPxHdFz+4mKylGAzzG5XJPO2QOv52RR+jx7iGiGZD2dw4uGiYFAimsvEXW4EEnvJDmpu
wd9eiXCYX59UL7YqO3j/KNunxf9z3vdFaTvcGIhPop9TPf/SzhOnQ/GfwBNhd7hK8J0BihmYHZRH
+nzvPGw0P6h3jcJQ6LGGJSGCtXxofKy2VyRzhwoRHwofwXJyY0P9z3i6HF7abgNXwTiuiM8Rdkgj
evyPjEAZ6ARinVyRckGvJ1fsDKFxnsChFkN+SHb+BNIXKcLztYB5qBlFHwvLuh/AHfkXdu9vAPrJ
TO9UFYhErjf6Sy3nHUIuMHWJr/Qn7tLW1zjnBOE/M26pSFlHoVyjOIin/NrOwUWv29tGdyTzCIjQ
KWYv/2GHz82spH9FUOEX1z7mPYXNc7JEf6xd5zCB+EyLWspE/Jg4blYDtFrhVyBmXaN1SF9z4jcv
v8IFLME8tNgXJATfc9zYDGOjD2JRZilFzhTlIdfhU5Vs5X+ZtjARV9ygHK8k96N1hr2cjpL8KrvI
JDrN4cpvFDfgZ62AX2Onh0Eb9uQGjcWqFzcak7DPsS/d2WVjrgmk+E/d4c6rdLuR06d4XLQ9UNmI
N/qjimP9t6cNP7pLAkvyBqMP8OUFbxMJ6+q+l+dOb0vZ2wnodxthaTHn9XLmJh0g8qdWCQ71hqR8
jyurhI05w/wVObgokKkIyiHBMTv94rbMXxTemQZtZ8XMz7mZVNALQ35VDa5psQfw9y2DYyiX9nkf
3TZSQV30CMWq0hNPtViqylFXoitPEHTfpepn5K9ceyqKDiS/T/DFs2hS0btah/RkG7yUmDlhdHK7
S4XP4/VRRPwtGrz88k1z9pH43f6LWHR+AA+t2qChXdO3MaBoFNv+4ixMwbT+UKRzCQV0W7iRBcEp
WjY6xMKMMb8rOkPZzuZglYYA/ztYDcUqe4LOjOrtkryBn+hIaAEv5ioA4khRvEBar9c8x0x2tkJx
PhLQIa1brPBXFUJBNzlGCc6zn+Vk7KfHG++5yUx1W5weiHDzBrDOyFHpuHXItcghm9PpsOU8C0GO
BN2Hg4CbFdgPTuSfhhA4CaE4hTOagXoWGpDpjfzDbgZ++ZZYEYrL5NqZBl34pyeApkh/OatlZJjK
QLuL7IOrJA/zgo3PRJyxooFuJdP/pRJT8W7I4DmVf8bLorxyH7Csa5eyn5ZWbivZqYC3v9By8rM8
BLWQFYXsYUGrAEclJ7xhXCAVv/19l58wcmXadtgxTA+1/jPZgT404kQsYkjji2sLQyy4rn2TvtIA
ZrO3PtHffloMnFQJNUNOmZ0OpOWAOBvffoIq2v18tAALaFV3k4ru1c6BEGhjbcR5QFQp3uzXb/7k
dd9Gpzy8iUEGchqe2s4eNpI1TTvbdvodvkNTP7AqAnlqq2rAcb+6QtSQgX3nG7/DilcjIoXBFYNJ
1x30lFCEYLArTpGFXKbHMUJaLhiij6sV7XocEpAo9OZn1umQS5bcLOHPa1woLwTK+UHQ8E1ECYuk
u5O0ALR9pKZcXURjtkoINNDYtafM0T3uy9s1UMkS0U/iDUFqOWvfPwub1d6xhwKS8ptPBXoy9AAS
op2t6JbX6IyY4Cr1/P3XQQ30BmKarv3yDb9tSch6Yd75kR8QdYvpQcYTtjsqOtS6X0JdhmCz4p5P
2VDB+ZjnMMwCDhAi+0KhK39SCu/27/s+7cWz6antrpSbEMs4Ke6zNfxxhevvikb4u0EDxP1XcbdQ
SmOnTOzwwzY8KuMgE+kB6HYHSbKjIdTddJE5xq5yTQ8HGBEEfA/PWElQzzQ9PKwXAiU+Fcu/SR0o
shwA5+jZS5VRdLY/2jAnft6NZfVmtaFVsdgOEFhtrWRvlb7e7Pi/AHqviMNR13trzY8SB3VRuq4y
5QnwnfcH1v6TXNdnsF8pdlLcNCMLnz9FXHnb9TUMzfdkKbdD8Guu602LALom5EX/DNq5qGD/NFSF
n+3dvYHns4OpIRa6+a8aGvBdb6OamWHefnjg2dUj0qjpCKjuEYBJ51DQVv/FdLolexnIjrDY96ih
9TtPcfilcXLojwDjB+bIhyf3JL/s+87NrHiRVEjkqZU1GZomL83iEb0Bi7kjPceXh7GsUAwlNguc
/VJlPGVC4T2EGHjuBsiVQBw+hU7yt+lCW1wRx+qgjkDxrLA/22lMyp4grGuawqTLZPn16M1fGwuM
ALxMiDz5UDNHzbUdEZPZYLj07XvMulZFgAXlCavUhlHeNlo4AH1/rMtroz3nlDV3ogwTNheGGWkz
j3mepJSkls/kPCpmiIRniNx+0rCQkZ1aftR2VJVNBo1RawZRw5x06Q5CQHjOgjnmDPZ1pADDoHzP
E/4oCjiiukQ+w1yrxf/ppeeWxS2Ws3cncWSwJ3LmjxlqsQvxhXlLjnQujmq9RXd3SKzb4W3BT/+7
t6W5lVQmlvAgCRNcW9XF19a2XhMmMswZdYV++3sQ8Xb11hOj3RbNAXQ7riiAEmiVp2F1q8ER5Zo8
YSZWUmn4ZpwGS7dFa45Jp5FEfdHfAL2s0Fh+I8NIaVfomVCEfcy5aYAYWNjuF1wPk/uPdFpUNS5p
ybjxU1DedOD3FCmX4HrbjzpwhECxeGKy9h2T0l0jA+109oVVg4D4a7WVoZekU9W7QaYnIGbEamxW
q6ukeavZCtHP1UGlxAL83CGtroU5/GlLtiJiw1nbIHVzzWe710968zvSkZXaBRJdIcT/mIcQev8j
fUcHGT2MPspfX2Qo2kMB3738ifheHkspfcB0dJKwZ+doNZCBuR1NE3E5xncfiJixLaOR2MOI+MF6
QvR1lC/Pb569/Oc9qqhaxY5X7xHrtVuWoo+wIPNs5YUxBcjK/0gOWc8yPApX9yMGQh9qj13uux9B
GAW3XJZrc/Z8DKQgxpO2A8Z8PNmTjiLhcZ9p5kChxDHo0GEBf3+m2iHEVxiJGxJk0HvXImjQ+/kz
dj4rcrxpwovVMi4d9dJB65qh3HZ0OUUTWSfPErJx0Qk/ke7aWuRA4iV/c3nZE45DfY2OTo43N1ex
NCfb0UxjidM1F52b2Rd9Qu2LA5bWWggUw9nVlpdvyVppCXdBp6GK6boR0Jcjm8kR4gFtUjtg/3x1
PomBzhLBcHRw/fIntCd/ARn1OMUyx+8V5KxWzMv5yOneSU5fDE1NvQS5Jo2tVII2Yy5ax99cciAe
3C5MP4/DAo0uWTBMgm4R48w2/8P/lfB/TgmG2TWtBmfiJsKbFuYBoEWFq+qmxFBDQ8SsnV6xqZBb
3htnaWfu57vLltpk7BU43djzr0COc0I0N4KVcX5mhmsB/h1y1djc6BESebZY3qtHX6qBw2IhMKF2
HMofn5fIDQvV/wmH19r6dacjBbTLHfsBAbkBOO3LH81o5CelZ3LYVKDNbwgY/Vbb87CNY1G53dhq
Ozqd4+jLvIhKbpONJNErm801X8zAkuuZlB4MbC3V+VFhIKSfA7UIGeWlf36pjUh8est9eMVVBrTI
1OsO+17lk+WhhKn8NCuM5vuEAyHvzGEFjpMEwVy6/xxkq0DBDzDRvPqhbXw2+U7RmUSt6E8a1iaJ
p63ifnZfxJ5E9wo9UsZK3Htd4B/B78Ac5d6wf4e9n5bGWA5bE8ra+E/uF0m1W+B1ZSBOsyF3xx5x
1OkplDf+knyjRTSwjobG1qjMKS543TsXAAeawbG6YpOAYmFj70xf0WU5kfm4mKX8dKgjaNf+rmEq
gep+Qa8bgAYwZ06PE4SqHPQGMLVEs6L+vioM/4mD99aLbVj0ezqD7Fiyy6zxx3CiEk1VRCGcbFu8
RQVO0IcYvJ8OtgD/1XlPqt3RP2VLyooo2vyy/kqdUKCDuRsfmINMsCfANUgICoEzRPxStV6R6875
gel7Z2wt5JpViCF9SfxhRGSA44fYqhUCjD6fIwWE7Xrkl1KWYoYv+cdBDZ5p6m7NJ6nahlKYCmS2
pVKFAxRV8ljGl6MgsCBz/EOmrjcaCfoJ+cc6Mr08zAFoKcI5VHvup1KIPfdTREuXU77n86RStVMy
mK0X7ZJGtMZdfaCMB9eLM9Fx2Rna5ul4yF7fvEYBhOCyklRyLtrYNub+f2B6xbtXOdtDSIY7gBrn
zWf9YcHolbDUhCTJkatO2nlWooNHLFZvaxv5cLdMDk0XcT5qVVjWVujyBjb2fz+gqPJiiQQ0fCgk
w9O2wEkoEn+Pxd5oqaXH+CC2ZrIckOsYdh/kZ6bN9L1Gk2EejdGlpfrSY1y8cYdTbkE2vUbQCvbp
Gx+qXTmFXM+X+B1KzOgN5LasQnVMfKrB6Fi66J8qe1C5/9b1zIxOWcF1eKYgaxOB53P5XRZJqwqI
4/p9ojGbCZSLwPZaZ0/hTx2HYfkyAKyZ/BtJ7TBZ3uEfaw0WNQMFJiUX97WUd4OjGJbWRgJwZJ3U
/7pPzi368jRluGqaNO+7f8xJ7V8A19qdUi88Z1Y507NjpmwyFNYy5ifpvBYtCYA+ixZGQ/CeFqCL
2OMPoFk/SKG0b1Q3/pEJXbkqqcSEA2IQ+dtdbyiLGCgQRxvV7zAly4A/9VazmV25b4w3ilSUFWnL
oyqMY7ySfVtH6qsdOQ12+vv1JUKpVtt2vIYyVMhHYgPAZ6O+kWn7DfBBCMDG6GV81XXE4rdojcWA
WEHUT8cTM6ZvhRq/6uXZDfuN9ULfobSH7/QGjhCL9iQLIdBkYHKU3i8Dqyp6W18jBWpv3tGf/O3l
JnCxeCXnggTE09DA9PJJXHV02tFS6xVIxzbMhvzwTM7MQLRCcsCd+DQDpUV9SNWJsX1F+DofCq6k
s1+96Ea6t13w54b9xMHkZUuFv96KFR+gv7UeJG5njQWzOnlmbwITnMClsywO+DpNlXKxUJiWSR6s
KYth/Ict5+25aaAEz663Czeh035y43aTmxSVvLSFHIRIw3VgJzK+f98BGjvVukQ4aldZtbOVvBEu
vl4LI9R8TjktFkm2MeTQH+INc+8B2QmJ1T7yqEgWYeDES71rVZOgxIU6NDtmRNnCXe4pzzBfwV7u
Noi0N7ptKkeBL5ko8qvgW9x99n9kRHiU/GcL3wA9oW7DFwe++0hFwCH1KUKokOsuAn2Hzk51ajQh
Ztp1PbiFxxV9uzy9RLrKEvN8GkhOcHni2f37gKIwc7cZNrKUa7/JkbgAWt2go39Ognf7vieLZf8+
PA4ff/mIkTy7GkzWkdzoPeRdvGKxXjX7VsP8G9A7VFl954sn+M/xrXWQ8LLhdwv4/UeBPPOnBRMV
LhXzhGu+8lKnRwcZBUD+WsYTUyuvGoqPdRMCTVJv85Ug+2kl0qzgyaQCI+Gytqkwce8xpyyMq2Ti
QUNLK+vW8w3fp84QydGKBcNpI+jzZgBpLWRFZmI0VqEiv0VfiIjIxVjOYKT93p5y1QRbGfPvEti9
ivPC7cYYApnctd7+8alPHWn3V4wLmycZbrSYpQBDE9XcZEiA9ZivM2OnLhuxEtyoESRBq8eU7jvn
Ka1iIcxzxPOjRYfDdUOjOeIEVkhG7+74MY41zhCqpuGI3JMr9OktQ9z+f3h+2139QtIcc+kJoUYW
7oB2AGMXx3n4yrkizIMDzGTO90DRcbc2QmGkbXQpbeo6aQslQejrGVx9Hf+6jUP83EyQIPNP7D1p
Cq6t1G/EkxqFeMJKrqKdURI9SiJBQXyF6kbHanw4L16wpU5tiD5jMU3svyBYDXxp0STEZjqWVyCW
XxTHVT2t3to/rjoRXfmkc4zBwCwmvbPdIgci1RqCzim/qXj9qmyG+D7evKW9JmCLi8x2VPNH7q2x
JMzVEAB9hQASJ67t1+E6hpi4Xv+I0KJ0Rk2/1l+8oqDGJP4gyjatzoU8ffqUsJZLQwJF8/j4mM/w
3khvu9owzuuCuAAioW9x3nc0qZsWFpXpTcV52QsRrHMeldppar4JWLijIijQewjpL7/JP8fAuD5i
/6fiRJv6KImKbixIJ9MFERoaoluptzTobK9Rc+VKiegB5xs8ilPxHdAgvxHb+GcYvmYEir153BQz
PiqHRClLRlrafjIyPrhh5m1lG0pRMD2G0I0Nk2mC2Ch341AWViraJtRn5c5ZTkJaogPlP/ivI6Pm
1QbGkoGzfrGLH9+b1HpWiel+HtN9DypsD9qEpFOVNDIV+QteHsEdePOuybKODMa0iNIdasJ7Y5E1
8ppTX9C8mC77A8Ub36v3C4rfj41sKKXfMGE9A99bCDOfE1dlqzvfjX+CkuLDhPULEpwlfvahVUAr
VOj7qmXU4B6/csoRAWO0EDFCqAS2MlCEKfAcxOrS0m3WDqHpPSL8lTD6YvjZ43ivCohTozBMRIy0
MBUkY/ScmKEh5WhQIgezNg9hjPNnugly+4NIrbB31NMSx5ctvG5LsGZ+NBpP+zmDdUFYrpg38Xcp
Qs6CN2WO1dTDfcbAWcEVytIDWBaK2bYQaqqByDJ7mqRgeZd40NSv6wJGo9fVhaRKnw8UTZZViSlc
89JGvny/x+QQRJnK5GTvimlSAtqOcwrjE+qm9FcQX/A4hAiwhp0WwUZ3aKdait6XRy4NIuvXi+hq
CUmupo98wt7X9aSB4fV1c10r7ZG5pV+CaaIjs9/pWUL7q79ID9tjCP4/iP53a5Qe+BevRiytWj0Q
xUOVyXY7F6tkLAJhHRVXNWRbfs7Z05kUpnT0gee0MZo2CEIO1dI5HrrhF7jiDspaj7ovVgK3yuMq
AstssRTk4x/8rVPuz/e1ZkE4t7mrdkR0YMWCuCq/SED9mBQIBtRZx/yuIAUHzGTAA9zByKb53MKg
IBCaGsyJObaQtiCN6b5DfrT7rPdei05F+BEIHfmVBG5F/7IsSqf4BTAP32jkJmZCMJs8mrAPF8Bu
g0umiQ+smvH6CkXwiGM9F4n11kPbRizBAmkSjLtc1A4IJYTmhFiXtBur1jLex4e1ztyBhx7qOUPi
WzjXfeNugglvlauQdE3CrClL9PoFrSo0fz8oFuK0nZnou2Qky2ntTtTFcbAeEuC96XD3Gp1bbGPl
qjbYwZLzW8WGwOvHtMPI62/dUMufSN3BUE7gFiCQqIuuc2TwfivdewKK3wZBEFAj7Jp8N0LOCzyc
oTskyXVo5UPbkfMBlUnW5F/xoc6Qwo8qYOYf5AH6Bs1biNWD5uylUGuLasHedcWug0GKjwJEBlLq
s7vXdJCzpflvX8wx3Nt8Jz3KhoDPTMxP6PSmS6/GG+t4utr0RUWdimCaOLboo/js3x9+kgOu5DuW
gCqTccFQwF/QGr6JP8bejufjzn2qLdN0sHftL1D9yobjjfh63r8EMPWclbxNVKGt5Fze1n7XotvZ
/btUYW2DbKXzD4RicTHkm1R0I1XAlVb1YejnbRA9BtuwFdEieML+gA51K0NMUfp7YKxtThLOddwh
7+SFRG4RVxJimSe9f0oiLRORLyOXqzGdBAtsalZHwPtFLAv0ZLD+ConV8Ma1nj25EsKhM/4UY8ZQ
euTe9HVeEP3YMT6SZsSkqoe1Ik7mliJ3oWpXOc8Ut8XFs8Lhxj9a5K9nnIQjbh5c+WxqMUxlGBhA
8qGnqb5rsiVCOY6EUkyX3o8FzaK8RN9d8vSI1ZFQkaYsE82+8DAoVPbSUFX5Saw1Rg24zNRmUz9J
w00jhAp8Z7H4c6rf2rkGn4WjAj4zLwksogSxUlVetgFzckpT4aZVWz2VQpsDyp2VrIsbbqLP48WJ
wmRv/Ip9i767a+ITiA6/8EaxVDmTGhywd41/9nKtlDXU/qaU/Q1Ak/ZP5L9dEGnEsXN7mEVauULQ
Rd+C7GZgI4Y4+SvrGw+aHFSPmGjuxTKzSolkfUw28xVW8iDWUL1w8r7soNjPqBIXS4nZSlsYSgTU
Z0uggEGIz/NmudRG8uVLLSXcNF7zr2+EGXEx7hPNk3QZHMifefyX536EE5tQT5+hzWMVoJw/6+OS
O/4Qx4W4ZlLzDG1HvRup8g3t8099wQdeeQeri5SklppXZzyiJb+GSaplqHKDX3zdsv5llLb9bUko
+njhHHRtpzOdi5kCK3yEhdZKqd2Hl61eFW0wPOHWkXMYqS2WM9a22nlLev/Usn3JpfatIsLdZ6Rc
nT38R3SecPhi7slWwSoouCjo//IU7Ocrr9+kwAFLEsi8jf8vJy4FPUcyCrvFR+ZCh/yCH/6tpi2d
/O5yhctCKqox/6keFtiCiMQzsph+aTf1F60Kgsnv31V961im9EcFTzVx9PL6CzQnBTrEOmgGOCvx
JTtcX5cVgbPAK7Vf5aAu9XTKVMECDya4PTDg1v6D42NNObjfW6FKf1ds8Va5qcpaclGnnfZdgTf1
5pWHmEhOxWjgQO8Du6kBcvAO5iTOX4z8ohd5I0s1A1M2bxQmrmCfVh5GpwNhHJGNOYqidiGCCX/h
ISVscIyuit5pzZEtUwcoNIMlWk9q67+IsxPISaM5TCqmJY+WyG5TPTKQnYbnVUSh/8/II72leVVN
7CS4YDfTd/eppMWRPjyLiOonGPQif5M5Pz4U8JiSwzvRAMAwEI4RPGF81PkVdWsz8tG7MAuVZU1p
NR1iNm/dZVCiAnXNaadiE/9p7EQLgdqGdFjyb/V9CEsy97OfLdpb7hbU12jbCG7blAsmPNvMrReD
DfjiFZs+IvPuQfal30JBgc/mDao+7oDwDNAmG0KnmDHL+z5jYaT1AEhBV8Ac8KYI+ITSRUO6VJZT
lwvUGtqBgmwuSnJWtGdU8C9vl7NlWEnZmGrStaZzSYvRVdNDS3T4aap+sKrRgGrlDnGagmPA7E0E
xQ9M9/cLieTDM/KU4nUzmm8QQvFnQgKQH+pUAZKyEhs5Ua+9EOdxKb9dI7R6BuZdpNMldp2YOxi8
U/+TY4dgppWujup7LNh5Q/ZyqzYLagq3bVFTsR6+YnAvighHt7eTnHPsXFD/G7fx/yT0rw7vbqVI
GS45o/6JqS+agMiQTlxqLYUKCCGQwAb/JxprZ9v6MpYwyMtCwtQc3ECY0nd2BRUSfMvZbVixbz03
x8ThpFkNSndsoZb2MxrPURE8ZU7GuBIO9m0EBk+XvfwOCkYYOUd9M4odSx3VunIHj6bN2XUk677V
Zj/TOP/n/Z7vd7vtUqXpp9QBUrsZNyrs7a0GRdZysIRMbgKscYIDBYK/bgVHtDEv25/S2ncHXlhe
S5GiTKzsomvHUz76xkhIF3gUkezwq1r/9Jl0exD7K3Nx8Z1mKFsWhPkpzCM7f8tkdNUnX3uuzLC2
wUp8TsONP3j9+Zxv7Hrv0AwwYSljwwhSKENlAnenretl1di/NasRN1Srl+2itBrJu0E8D+aDQVuv
LQk4viOR8SjsO6wda9rHr3Op6ydg2oRU5vWPi402n/PA9slRyilkqur7RxwYsj+1DWSpUiKqiSYC
fGzutyrf6O9PZT1S29yaiiFa5UZfsHrHjKoo8vWaKlByWFYFhiiZV0vLYnKkLT0WV2RqCnj2fYS9
XA+a2AsFQM4Q3snrsLu0b+b4KcpXjgcCX0p6MLbZ2i9/WzvExunzQ2YoNWlaeFjhNNMlJ3EUC2g/
Fe0a4YZ5G0S/owYKhigmvRu2ouNfe4cHIcAx2P0p1HW9LxNf5/Mssb4viM773v4lxb4g4TwC1Q0y
7kwbldA4Kl1pkvM1JyBo1QXJhD/qNNpbpqLFfX6FnXzjfihIrlGRwHiVQI8eHrnKe5iuuSBcDJLB
ud4sF0GOdNNmpAeslnYPnYtH5m7qxxVZIBYGjZKWbCbKFdOPuGzjB4xddC7ExYMdQbDFJrt1Lssm
r20NjGSxbQHMVFub3WsSgPvrCT78trf/kwFwjq4dtJS6z6XfPC8qRO04HCRRctmZ2zet8ilT6biR
YJVNyz6l6NnV2YztrcCtDC2/d2uFn3KpkIQUzykJFt20za2nDl1p8SNWS/r0Md5wDDM1KVeZoN8u
pEM8ZCNTb+a7a5IKVKqZRmUB8PgnJlM7gjCVMy0fIxy4nkck73CfZ/gclUyHzdLHJkCO+hfNMLLl
T+S/pa8SA2Xfvp/a0J17YU/wuElIlw4ABaQU0klrNURQ2dHDK0atu+Z1WWf11VjaiMZMVQy8EgNf
ennX6V/CY7BPqQO96EN16znnePSm1aS2BTFmlnoZWNYJDb2Ak3X/NlS3l3JmPxShzNbZwuTdC70z
y+MySbEWWEDRU0oNNDmYfY3tW+VlXnqLbwxe05bqoGQ8lWYutKeFQuAXTNSUTKt/i9tbu0QCD7g/
LyqnT5uVR27BtwD+gAR+I3GrCN2AwLYKgTZYLCcldsWbVSh0tjVUzHIrX4yCRjBXElWFZPsXHWA2
flhMQlfK7w3qh78F4hpxpdXDnst7ih7JNxXmFpsHdyBoPYz5hEd3N1FCMTwn3COoWF3AMrs0wbpk
5vd+hdZypLLkdXUcJGmWdP0K+FnEx2YCBdaz2xNgTgPGgiIv4fKb150gVbgH2rE458Llp8Jit0+a
CK2R+0/DyKolPW9QEJ9ZH4RciEHZ6fwKlM7HuPR3QYIGyDhKHmlX8CNFnGCnvP+l3KPD339224Hk
X11sdO5Zb2XG1cAq6T3ijztuJh+hZjJi4CnDx2MoToW145+p8jU4oxWAb19ZiKza20ACzVUBJ9VB
7G23e828I6Crp+H+EloIFzXpepHhiiXNDZEr54yQfG3UX+Ym/T7QOR8YBqlcsNWMLfhE3qbnrxtM
qVtYTxqc9QVUcy/j/CUzqTDiVi5z4R9eLG6xdnV56910bCJf0WoH/tgaqsTTSsh7efrF16Hm7Swu
ZvKAIZ6hJDI1RqxUAs3WVFB82hbIfX5cI7Q2SJId4vm3l6hwVX78B3jQQs7cO6sD2OWn9PxqD4BF
6k+5C08lKXaHl8eGVet0T4uO09+CO7v341G2uB65mCLPmn4w4mCTcP4jxkvRaiZ8NOsNYR05FjH9
16HLvK1g9kq9DmmLSBqxvSnJ8kuVMXh8xg7oWdfyRtLOIto2ffeVgGymAmX+s/uoDGq/WO2m/OPq
y1Wd8uZbeuInGKRQppLNh3QExhYcCGA15o7qzin8CCvgUaLl1H00g88H2eedllpJwb895F7wD8DG
q9l3GW72h7Pt+aiPODSrxRJ13qly3oowVF6OcjYt/gk7zOvtZcqKyGogUbCKxaD9+OjkKoeYe5n3
qTEFg14wXMXTlSGqnEG3vvzYajMCn6fZU0JAI3P1EoYgfjVbUApYW2y5KiWEaz0l8CX2H2p2VvU8
duOYuT5dPNcQL/MFxXy2/QnUYjupIXMEECOIRSPQ4LqVOA0RmT0GSiWMKOrE4HLrGyX3jWx3G8zH
OXPGyIXpSMfmDj9OjTm3Wo2xvb8dvl1R40Y3zjMKY5c4MvSVVLrQAqu6vlOLPMwVV2PWnhgL+V57
wgoGI4vF7T6rEDcv2NjoF5VURS2881ZtUZ26l4SkWx29uhLqDiQIs70MPfpcOp4VlXPV0oLVnuh9
WwOrjJ4o+lOGmM3IkeZMjG7OpCyEz0LCVqc5GsyXRiqfeBC1dqy43lw17y+FoWTKYulhznu567FH
4NILMR1atHTE2vnYtYYvLLmyOce9Qo/9jIqS98g7ol8Z+KUKyDyeZ4OjWnsOG+COUlmRJ6uM7dgg
VbWJ5fHupuLdFD3Seauqtsjhn+rpICRPYKZ+MSvqvFC723/8bbT80bIw/mAP1trBLPYqo5fMFxoi
zrDYjorWTcwynlYYwZ05ccoA10O1URW2SuByu+Gx8kkY2DswOEi+OQmsrWpXk4WtBxU2uquZrxHT
J9WjGG6PSunPF1iBSrj8pAQAIrvs7H2sHzSy+gjUNB9Vwp1OQZ6c8BJ/lfAhvIFbH5xUNk8EAxMI
Dp6WbfQ5qY7CR5DkiDRlr7Y193XHZWROSZWbM2SE23MYZQu8iyhWs5E0CnkCkJIFoqTV/5c6nxZ8
hq1pqOnUrxCXEbUy/qN9v1mW+DypAygmGwfgAHWythL9efdULQ7J/m1/nYqucLT3DDzLFsC+li+G
3COZK/7fkQirXh5aGF3+nmGki8N4Dlxb/noHODl6g9xFxq/xsLRUnZjarO3RuIFpoMjJGod8G8gq
izh6MvWW5GybR2aILv+SvuN2a6LKrMPkqIhf1spM2mFmAt/2MJBY7wvYyTI5bfniKnEx3eN5IcOZ
zT4VF4fzOdOwAR91ihXXcjWW+VIhWP5YlkmxyFaviMAeFIqOSS6gThT+tCppDffF1/I2+ZA9f8hp
xV5hy4RdrYACNfmZpmLfmrczpP+CChhOKd/fUoMdEF3YkDGglwk0Zwc4fu3i9lOigZ/ropzWzglU
DOIUA1NUYQFoyqejMVrqPh79F2w7Bi0ZPRKzeS/gPZYGxcNsbBKxu0FJJZk4L+Vx1V003eDWGqUr
Qk2at8E6/iTuPxN1myrJWKRVfQ47Fp6LmaPjJ5t5uwp8r1IycQ+MUPFRtT1t6SdGlDQqGtQ9Aj00
ftUwuQUJ/FPbvPKd+b7lIOveT47GxgOP12zdo0d5GVTeBxgkRxOV2jWRrefOswufHQ8RzpQy+GBd
o9YXpuF6YdbN7vIHrLP9cSvHHe+jPnI04ggGrAgqnZJp6GuFrrEY7rdstIPFrJegNcpGE0RpmbYH
zMnmu6YBAUf7U3aw54UZjAAbQ2MtL03NPc61PAMqyP/q+ufeSeTkTDD0YcADDz1tkei69HpPQy9O
UuVdXFGCF59CVbWOzaWvb0W4329yx1sgn7vZ7WDhQinmksDSC1A+PWvwyp7Vuuj/VyZA7hgYJ5aT
09QHV0ZyDA5x4BkyGy32fcnzVkZDGL+tE1PnUUCEn6Fg0iC04nbFKc7+6CJOpe5mgQ08gYxgHh7R
YVdZVJ7FIEHGsITM/cwc2nkr1TZ3RlVeuw3/rGOR/267qnUUOGAsJk07TPhJx8LP5ZEJli+hU2ro
I/XIz0SxFo1tLgOtSTc335MYNGrZD16XJNY7XDeCWTjISAz0ZZvNYwXbKIUKCceFQ1vU4mKWLe0Z
mHVuoyqvpc7uSTgxcbr2KaKtauvtFHQGMyih6IT/1Ccz4daRv3sjTpb1sBAdgyuo2NqaLhH/cVuT
HQFGKBhUTlRM/6fTcqIU6JroxBOK6i7sYMnWT8tgY6UZ4zWX8yfI54qdAkwJzUJnq9k9RGY/SAcm
w7rQ+qumQt7khRBcPY88fLn3E/QAyS8OA4hxOVSkt1rqgoNgDjxlOcfqrI398nocsuShkWDFbVAF
CaDPnmaNnEInwfLslOwDgIHEC4E2OCudENgG9bjr5QsP4NWcIcWE/cBIKg5Z2WZenI1zT8jas12v
6auoCsvVkT9R2piOOcUqGd4DR/Klq/ByMWvEglABNEeH34Kp23A9pvl/8sxdgVfzr6XJwMTVg5EN
Z53kfKKDk/0sx6beI/nfglP8L6CHg7bK/qT9+z6vNpAle1MUiTvSpD7o6ivvdwijFl016VTvXoVs
209+6Q9oNSOLP/6UrnkC02PTpUjZ+iHLu5qW4RPx3cgVOpKDp9NThbKYPVN7MZM/phTtuofs6wNq
zByz5Wjwi/P39sgMk3Xyd6waAZQV56F184lA5VlWl3gitCUjw64+AuGMdPImZZHkBc10zwK3XdgQ
bovnn6SY4300Ibl6SK8PR33oplyji5N08+n0ect6oUn3/3cZUGAn3ZSNLpol6i6DGZW/DwfXH+KF
1fcilADF9yfsX0UeGjHzyD/4x2Z2cgCgOrMa9SicwF13d771zfCOXELlFcFn/WS5fm29kMlaABPA
ru6x/s7h2VTrJD+RFlhLzaQ5W2MlUsPutB0OYczpzfXKZGMzoRGu6pBWrfNPu4+R5k6fJ9tyaFqz
SE63bPY2flagWsAG7g3IuqXtbBVjQpoY+v8LiGWPgmTp68grwQq6EclJ4IIRogVAlU5syX8mbxFW
PRMAH5zKXPSx54TxK8mcTX46wWqjUFEUMrwRVO2ZKT3xqqRYj9VGv0mdcEKiCshTSCi8044z01zi
L3ykEuSmeB/J/ZFvzmEJ9ix2tK1XsOu8optaYyTnHIxPuhlkPhG9sOOYyWSanZMObW7BAsRsGDuW
KRSP/HgU1Oy8+0LnTaOsnF5gq0D/uKq3TeWtnTON16h6lGcC8AHtND5urZcjUde+vBuVkgl/kgs7
vpxmzDz9aVD2gmtLYXFh94d1xmJdqo1koYcd4ILKYhx0qfPzWjrs8LzU4QVQBEwL+0xesoH+Ipw6
M8ysOBIov2f1rOcUDrt5c4b4cNJXnhc53M78N9t3M9qv3zArIdqr/6dEGy7nWcfsoecTyZADdv4w
aHHvJ9LYNCjsjCWlrbqvuwBe7HTd8WjVimSCXzl8SDLcKl1A6VcRPcpeB719Q9OA8zb9X8E68IF8
9yuTPdQ0OXheAIIXziFRj6ninmnF5FM9xQOc1zf4nvdTtD5VGOiKPRjMz59B7Cipb+cgOxgO3Z+j
SW6ECg/2Daba2iLFtd42I5An86FL8zASxdHpoouagAddqxzeJ09ZfptUk2qQugUaWjiZ6VlK21Wd
uLE1OnloExvg80qia+rUQoyO6le1M1qbsuONSQnW43ycOCWopGiMOXqO0GmyvtyjQFCd1uBPCszf
fWznTbzOe6+S+ntCuQdTdfoxJaIHM9FCxoFpTpQLlBzkrIQwzizCJTvCTNcIf9j1HS9CQ0QeH5An
ogODyVkxofskZ+uLBHOSgnIcCr/wS8j6xYrN/CXMsYABPiF/0PNfP5n3EWR/YNwaXqnCOuBUKIrs
O2oGFFvmtmgmCotKMGdPS/ERflQhc1MXz5Ulf+AKvRjy3kxFmy5klc7Y3UgJjW5Rb9PCpFzO9IAc
dS8d5GSCST1CiImzWWPH2P06LhqY7aGyAiUH/UEqUuC9/fIs0TtrCpoWXDbk8oPMJBNHoEEAsQ2G
g0OgW2gYDrOe1gVQUIuAeL1M8z7aDzJ1VIf9Yz7icLRtGmfR+ENBIA7e4/LoPc5fxiVY6WRjLh1v
QzbsdWjWcVXbwt72QinkgTepiVvr1j6EaICPCVc/B+e5ypCdNmFEpjpFwOwDSuJwk+gmLkVncwF2
lkZqPr9p1lN7+1ZFLJaPVjs5ZfZyOB4XeeNalKrtbUd0Efn2KIdd8k+M+YgqVwSwl4EfVqfTlquN
bz6umz9nnifVeLP5gOSifjpwcLPpRxZ6jr0ZBh6jq2ihD8gaBbe7/Pn0OXrmAJEn6QRYvJ9Ck5hC
ZFs7/gXz8JCKnUgN/KyIlVW7zI2xPopWuhXq9Hjx7rwNnUYt2CQwlV3Xf8jiS93a7OxpHxqI46is
6BG7diHnTCbzWIWK8xKWgGLVY/TBAYlnlhc7AP4ZND/fThohD9n2VEfUvWsP4xixxlSipc+ORqDJ
TkimRFCKSjtnwfHgrYqMPuR6yWX8DQ27VTvGSfLoipndFOvKDAI6AomdF+5xJE1tj7NU0klq+Iy2
U0t6hPMiZQ1Bc9bc5ajoiNnz+aYdMFm3T7ih0ef6hPKDNmlabtHzie/1bb5xToUj2pKSLDmf7M60
izuPiLdiiQl02npSMFM3H0f3j6kcmCUCb8/McuBeP4v926n20aInIKQyB6gC+LnYaOF6nQhFPTgw
sdPuPPWLCzPF14lKISlsCfazaIaM9tEFX9AkuTryOM72pyi+iyKcN+tqjl9kuueYd8uahXT79Fev
A2w178wGdendoxDzE/LJl4FCNWCs1ilYxOop4ZWxA+J8gfmqHSJPqwmOtXu/LG402mDqSBcKDakD
6L4kpVFtugyh83hUkBrt2T0u+cdxBSWZq0+yDE6dNFACPXTM5rbNPP+DdWsjm6zeWVyMTGjDFM6I
VjwD8Es2lurMsRcBlELRlmNT+DnRyor0RmfrvJ2PYbXv5GqXJrV7XSxvYt2bLvMoyOte9l7L7h3C
NzaCobzUM2J6LYkUkzvJuc1ZzB9I6ytyiX+cmSCp6QJ93IHTdjdFxme09kCTdUcWnvDSnOKxyBf9
TOXi8GbwNsmLjw53vVSZiQj2b7qQi2lrCc8dl7ySU7E+W7WI0Q9Jm4ei0o0H17iHvQp8FqGWl+VD
9D2ro6vJl5WF1wwrN471SmmryHxBlS954E6nL2cCwVSdAlu0XuBSuFKxQDrSDIzOspKPTkR4CrzI
VPpw1OYeaMuwclX170T5J/e7Kx3XAMrv7YodlPlqfc9hllU9k9VymRaxjptt4FYwsqSIBa7LGsrX
KkhLCe1AmXtz7/QRY67pkeWwfIXfI9luA97snmqE84v7T7+AbpMsgDDBqKbLnl+ri9CPVWeLgs7z
YB8yupAph7XY9CySs1aqQ/f1SkA845bC4jlxw1LFevDhS1PsAq2CRib/eAqeMzY1AVmXc1WdhbN0
uzBbE5Z4XhqyTIWdx6/k+/rLhrudCgxCldUQAa98XCXT7vDJTqP58+l8LGEZ1/RqVy0BmKu2Bpt0
iUePaAjFUGppjKlOo/0RQCQV5BcH7d8IGL4jb48WXp1vnrqgljlYVA1cjEeUoswLkBob8fxcNsWN
FmR52O96Y3wBJyr6BCdR5vNFCmTZNBIonRVPA1yAX2NahfyKHoMhVKNDNjCZYQfAZMK4Zqey8aUw
guIrEezH0UYtd1PbtW+0V9QqS4TN+8z4fnICcQXYPJW1lfMpyHBGu7ij6TeZCH7iZzcp+BSTfdQ5
nXJOGeHzqgEDFpXZFbN1obYEnKRFkWOLElijikOJbNGqkbNgXD07DAynZbRw3KFu/1IYYaIglbj0
/4qNffcTC1QwTnsWnYO1y/o+GJsF2xzWi0VIliQWJNRsV6jV/Py30OX04Eud//aaVUvBwMLtDWsa
kGmyaf1jjuBlahVT51q6zBgGbM/bEuNlY9S/ALna/XALfg6REAy+JnOFfJrCjSO+kui6cJx/lwW/
WaOBriCfxqrNhyMm3kAEBHU87PUXYB6gJ6eYgDjzAysh07xJUcSfkDmptjrazwAavIvq9rG3cArW
ucbxsRE/8DTcTOTi99OblgTz9nH/l+irxvjIlK7gEoiJLGZfbCV/jz5xpzw5TTBM+sU5MMGMpgUu
LcTnhNeuNEkFYSMn/Cc6qA6GUvau09JRYmtsqRaqD/4KpJOSIMox8vBwv6PVzxRDEr5JoQGJJHie
y50Lvn0IE0R45sjI2fgkmPLW3OTcj/V/oHbxZOfimoYD1r4ef/jGLoUMaYi3k1D7aAcwHzmnldsy
WjUMZO+hrkn6hnvnB51O6NyWlIuomo069MAPcYd+yAJlB67HT8HgzrJzrxkdNzBPAyKBOzbJ9PzZ
YM6riApwtJt6auTDhGvN931378vZTquSRtZGKEtvNPGQFeFFMYBuMKjPw+aUVM+i0bfFAvJwNpGv
5bVtZEGeSww+Kx9UnApNtoaO5hI2nHigCQX2RdcRznQ/1fYsGOABeTip6D3KxnGhzRieba11RzzF
msSvVWXr1fcQrmPSEQaLBMNoLNdEih0fTwI4PM2Z6gCl9vjqb/XQ9c5uj0m/MNISM1evcJJC5ePY
3oaq5E5Nt4SMjp1tFn8GDFZmUKmvG5834KjVniyobXF8hsCSK9545l8FYHfOpIKU2FIXr6ZC4cFW
6S+eaVl3EgDr56vGSeGi3jmpwRRcwxmgvEGsTKMfO2KSGbfOpxemB62Llm04rPRdmZUAQDlsIkO/
uIEuqVqOHJxejozSuhUQe7wBtx8GVrjwi8BZtMUxaDkmQBErX+PUAlbQ0nRi/yW6p3ZtdMIozsTI
rZAXcRVEpacemQYQf9/iHCj7Yuz1X6bNtezpNp3bBFwOO3uAwuU64rrpQYBmDOhkOkjXX0PYjjlr
03hpPXNcBPk2aLK9w0RcIaVfN/7C+fSHcZtncUSTApIQH9IWmFPKHP0K4NvvaCf5zJezlVEzhzdS
KcgD9mvAnkll5JjAzWT3whD1taiCJJ/Qlodhrns3MfpLVIXOtOyOoztlddtfSomQLsdBfd0gWOVM
s4YPH0wODxmC13ONlRXYZP1zAQiGQcu6gNrjVcNSjfh9Cenda9htfBsUEWH98nQUd+Bsw+jUu9NH
8ExYMZvCrRizNKHjvjvOQgN39hFZogh1d+yZAi34pb+l34DlpSadqaZ9PfpnEdBiPFZMtKsTpkxl
xuItZIHaLfjV5lPAe5Yn7SZCrVIOj5WKteXSBjEx9ZSY1XTUjOPBF+eh/1A/PPKSbBJQGGNJd+OY
5B16wLIWvCrSnICVAcF/WNWi0yCbHUeDmzvloo7tJFOA1wpDU7lEu2drvvXkYyRbcCLT6dJC6Cms
P5ruXlPnBeC1q2Qsh4fxapGPfsXWpX/tsdr+WTdGGGzCPnMritCEB9ZzmILZvNqSsuy8hFPhZALc
BKsjxqPTRiuPLUmENd1x3EfYFtXED1b71fQYC+eXuRXKmO20yd2KiAtPEtxkpeyzp1/xyubONSBn
WgSSaPcNlKeEI65QVL0II/01t2WggHVVQpwXvPrA6NF/mjBnD2ZgM080rbGITtURK62DJVpbAYZg
72qnFUqlfoQd7xqjMAYOuMna2rWIpJcH8enUMb03ItfNuH/CK/VBBE2uSyxw+vVXnwfAG1KAlVUb
rNWVFl71TQIPvtDZbnWwFre5VrixROPn3GF/nfM5ugXPBEwZBuWsPSsCGnc5VXR0Mp7Zj1eaAX/t
vYsZmrubf6ZyC7q2MX7flbPZbjPbAM0YT1gES4M36c60cjSmkO3628Rz7/NYuUVTfkvHG8wUN65g
lsXO3szycKVcnFCCdXs42ei34hvRMreKadWPz68/OjMxc4+b1Fd8oyrXgz9FgJtQ6Qj2mX+ggqcx
eHGAMTqCFlzAbBhTmVoePdZYOmuGVjJxxrnDifffuKSesn13i0gccsL93fF6rz3bbhNWoLJHNKys
ROWg/DKZmG46tP1TQz8rWwlbf3WgrPVNy9wnJfdqjUe2VlbykXes0TrGIyhh79grjggF2K6uVMgf
QVEZqzg9e9/mKwWZhtwM4E3paVDuut+Q3BLlfWPmEaIav/ibTWcFZK1f9B+iU6kBNQj0ohkwHcw1
T2cFZdQb9nDVUviILfnicxs/hp1r5iIC4oTrd42pc2BNFw7kCcQM5Bx1OqFZeAu9FFmx0z9RBrST
64n8vw2ImPbDJtfC0BT4sxClcesWJbXjGIW2CbkBI5FpPNkZbxajtEIoTrW3pFGaZNKP+LAMvVQD
0PxfuEUepmVhsxUG20r7QXgvtDB2YWuSSPgAJE30zImuYqC3oeiKMfeOF6OhFcaGGWtCHs5uz062
gtSWtVa6dz8ZjdCMF740TZtXlpiEPu4YNJXS0qafwTxvU7+6A2EEoB4J/KRLV6lZeVvVWDUMIMRz
y34+Ql1NaWydJ8JtpYMK/u4nE0aN/F6VSZ2H6S24w3GK9hc8CrvqxxgZv5341gIixvIDDEmKKVOW
SucDac9Jvp51V+xf4g4BG1LzKdXn/4+xDSDzv3f85StLYjo4+LJoDZT2oFBsmATDzuTXLV8I/kZw
HvW59w+EoVAwH6beCfdaDIoxS6AAgTApaQb4DZJvYI0NoS769YBLPVfDGoadv3OAiiTWavWbjX1b
ErKMrrdgAo+wbOlhJxkwCvzZFPEi/pOeDNRZrtG2ZTTPKEu28AFc42HIYlYnAoW5AUyjs/oUm1Ws
eJI6I/kx5KJ2V8osIucCx+TorYAjE3ZGxAT8LD6dpdoilXwD3KtKzYE2pBvqkFDvYHU7kb8wK2/J
033M1Noj4koDC26bL2KV/+duHYfOXmiG+9+MPXS9KhLA3DFtU4LNTOtywEnMhb16C+Q79YsETQuY
aiKXE4W5dmT9nByaAj9Lwh+avLm6ZVUJpR+82v+1EE1KzEp3GL6CJ5hu/6fnRu+FXlEB58snu+Y/
tybahqpAf08nbtUhnwwZdYdzl5QKudZOyAmbmL5T1VXNgrtEE700Mmkp/ljsgcsXE3G/9t+rmObQ
PvjVxcdjGctMV0bg5XTvSPkoUa1FwubNZDySht8fCFN0ndt3BlZXR05qjn17xXDaQ6Q3YWtX/1Qx
Qsuyj5yGnKd3VG27svmgvC/zlSKudjV7FdzEzCR7JlFnoh4+v8Y3ovBACBkwxteopx3rDQya9BsE
f2Laq//hgl252yxU3f0h1FB/99fnQvLryObmpW0Js4au084tcX6vDniaKCm4+IvgGrdP65pgPOO2
HzSCw4NDftWV7QmQm03GF1acRkMzqcJ2rtDABy1U2TYZ51hcfcHJSFIjD4YOdjTIVLKOpvJYGrwc
+URy0vmEku1Rj8tSM4tH5ueGs//3l/SoLmkjVcsHg5fhCr+TmrWydTeYWIhr4x/McdIbhUN7E6AH
sEMFgKOeqR5IW1vfF/gTNHWPu49BZqa5DbtqLJsZFqWN3S+1QO8c9WgfPmdHGkbaWBLXKqdug9Pb
+hwwDzo/qDWGAAsTv+tPPKlPZAXMStd3mbDEz2BTuvRATiM0nARaHfCpoxP4xodcKTyC0qjk6gxu
DKF1TgHOBozKx0vX+Mo7XDq3KtD2jNztsvHSisInT/MymQFHGVs4i651A91yoCihIT9+0FpA2CBv
BUt1OghJ057emz7qDnG0r5XEzyHphHokWda4W5gEzlhUM6Wjua/A7ymyijLy2YGnrTHruykNReVt
ftHDPGhwB7LAhubCRh716Dm1dgwNWzeep8i9Nl3rO2ntv+DaA4FCsIGocDlYaKFikuhlHW8kQ80w
Q3twNnqFaNEoetK2/PljEyyUoTt0aE/ANxBoMwMFG2OkuiYMszxNzJ5aeQ4BwXebU5iNpDrfeUmN
SvErPo2W1Pz1M57RpyQ8n1PxyxEJW5t5LYrBlyhdbU1iA30i9cVC2ceFr/Z5U/fPyO1G8CkacKAC
ozljgAItauVsVHz2ACMnaHSoZQHD0EuKEqJRYSqKqHgEf1l7qbx44galzwvp5gBRsd4DYaASdaYR
xytrH9s5L8SZ8N69kuRTJayLcJd6vNrzLuBiK2UlPzfNREfaB2h5G4+KjyHAMmuvbRyxsCUrkhmH
8ifsxImmCUuX2bxzB5dZztlvMuHXzA1xuzVs0xhtHIgLZ2O/eWsI0rdXWRPAEmMVQSa6VefiGfy9
dbNXRv2oDwAkjj/TBZl/4msyWgPu6+KAWM0yeqpZMi1aAa2nomO5ooVPqJ9ykUv13aaoAvmhjFqS
eHUwH0KBpbEQDvkRVo7WWKtCE1MEz1f83gj6XmJH35AQowRw0G40Hct6DPQ7CbOp7x7B45SPiE/7
l2RjskEGkitZc09DpT4MU9ofdSWUR1Qx2wVFd+HDdDVmP1eFlrRDmJa95GTh2EWtUL9j5+mQhTzl
VsNN6bZtU0np7xbwrYKDWwo9oVR49XbzUG/EYMw9ItLNXgjPyrFfoWFBLc4lCOaOvngDc6v+7Xt/
SqwVBG7Eu1NZjm/AfLgGQgUdJU4bZlfKUSs2dmulhZob7kPzy1zR/bqLqTM2tm7y905XLsqgOrdl
AIoPGq9pAtLjpqUafuNVOK0PfJcAN+OaF50u8OOANh/ptYzW3wTD2nbl999kxMPF3oXCRItFsxdN
qJkMZlAKMWC6Hms8Ee6QdH42HVmmaRUWO4EwkfXGrdhzcqxBLCO8Kp+2mceob0Zyv7DuwLRoNamz
IMoZQxZCb4aA42no3p6OmRBSl6gdKi//B2lqw0I0REj65/wWPbTryVHahy8w+3b/ojR8JZ3lJr/9
l3Ikw9mNP9VwG2GHvQGwSiNbTaX2f6lLMSxJjO3HsqMnwTEeI7G3Zz63C3hgL5/VtRtGQ/GUfBl1
v7bC/aoZtHR94DAx8wApVoq92ddMlCBA5CijGy3Htg2J4xixe6XcWOvNB9xFCIA8WKPcEmLwRD1k
6sReYrNYYIMIKwspXXoFC/5CRl4Me/PS1SG3ssHzSJRkUjnfs9OaB75ncN54myuGt+EQorSpZXmJ
S7q9WqTk107QXX4E9db9njRbA9EkhBXMttnxr8ngUqfupGdTeW/01PPSvpVjJpaoh2pVYwxinon5
zkhL2E0oem8KeAZ1jfWxBfdlE5vIUV/TQQwGiPaEHb7iSWxmViSTyT79bioAsoHyLurpZ2g0wZUF
D05Zn6QmTy0X32bNRyheAK+K+PRnasNnJ1eO27cI6niMMWIswa4iBiWWjqKR+D7N/8lI8mQstBbL
gudxuGvKlDhRToIqCgN6619YUbbhqHJqqFw4/YnqTKy5EaDhAcEPtuKboFz1Q7JLROxKXgL+Yt29
Ddm9xjJeyjXQYGswcqloI/NwzUwRVXpcWakHXJBPPUabd3M6kwuXZJOxkXhrUxTjJpgr+DL48/EO
1DfzQRvb79gsNpA0GC0UAbXnIMhkx7aqtZFknP/tsnmAk/CMoQRwcITLA4qSts7eCgQO4xT7h7W8
Zr14PeBhS02nKeJY+nd37cZe/cNpJiFG+Tvc6Jr3SGUGh1CCd/bWNF5fQjzS1/JrlUs2ZF+/E5Oj
QvfwDZXwtIa7tZEMKH6iSOrgVeF8qzjUBZXC1JprgfgdTveMRVZX1hHeScXJWk6DDEyUA2dWEazb
L4bK1OaUXrdiYk2T3c4xV/awB6EL264oU8EmxC1CzQ6Njsu5A2+EwHEhdXgqdLMfWJ+4C7z2I34Y
OmMVMdAMDjWP37/40kB+z/VSCM3qpeJnjVVV76jSQDxwXzek7nViF+onGFb7gCilqmefmAH9mxY9
P+myUqszZCfMRLTCfL5R+Zyiu00YKhWIJpEVv49hFfZ/tMVCxKj++bDa2EGu05U3fxw3EiRCguIT
ds/OPHcqN538dKNRgWrb4TSqWez2C0yyum0x46TAI8K8eYWVc5MBjmGzpVP6tBnw+2H6DYHMhbK1
T31orFi87EbY8UYn/u34pNEtWNRw9uzbCrj66EkdLV1p9Kr2DBK28m0zALbzgez8vIetA4y6Ftyb
adarIbga2+sRjmESRjlW1YGrRamcz/EfnWB2FzEPkUMAmbyznyui/LAMyudUkPbt4RGRIh/Y7z0b
NsaoIg2GuDArLpBxHjnIvN0SDPTc3LIPh3fM8XciIa5BMtvIv1vrRkFvMVTRtTeDtb9YizpYChrx
em7fSm4r6L5lnmZ/0COcb+BXJAa6fcG+jEAQyQwS5nsU3/kPNR2CHPKqrT9eT2WlZCR3vmDXHP3v
7hm0CA5j73YFmRJriT98P7moLJa0qptII3r3dcUNqEDRrHzDsK8NIoylxlM13n8B/M1zMQs/TZmT
g3QNv72SMAVFv2lOOEqrZFOyGu57q/PztL+WkQpQqclMZLYPWVzYnNR424PrdIBsEwttbb5kDZTU
wbPhnWgCcf3lxNPrurPxZwYEF1EP8ssu0EFiR9/gr+Onabs/jdYJrHp5tirSeKYNXX1D3OWoOaDA
N78y02uvABECi87lW+4v0n5PqazkX2gfWkvcjXIYNS9s4F0PKcvZmdNU22IJQQWt7Wkxcmnbmw8A
1Wy/cJGeGS1e9Sc3nANw1Jk/9KLMdXc5AINDooMRAm4fbHX2QilNJ7ywkK9qEvPyzQhYrA3dKzcy
Lh7/heh/i3UOpsImw7uo/UlorLKMctAPkz6pTfNGQKtYRaNfQjltEqZTlsTEjU0NaDShsWbisgBH
RDG21775Pqrv8txAGKZ4okq6Y4Dt7HyomdB2dcbw8lGjPHjefQYs+Bk3p/yvkmN3gm3KeBD2NP2U
c6mgptRDBMNDPV3dgSpGSLWNxnH+MISuVUvVamUb2ZskxoKf5V5hkUOUUzkM81ZCYtj5niDKlhJM
0ZjvLjQhBq672IJHO29Z83ZhChP8jGsDK4QoAycM8NuO5bIjS0wQv5A1QpdARdnjSXxdz4JpgA9D
XfxBhw0T68KOqHVY6n+i79Vojq5c4F54eJsvwVDeWWmHefK4p3bjPQUV1OZKcH8rqTuhnbiFTW04
MG7vYiUYj1ikNcTL49B5QpqRy11JjhtpB8Ga1OwJiCqrKzaUIN3VfSHLV9O5m0hYtXkqoLeEbypU
/iAqqNV6yra2V17Io9DM5n+sI31GOyL6wgikj2jbu9XHsaRl413Xi7CyK2bPFw1QAORcbLEL6Gab
nT4ZV1o/ZSY2ubsk+0SttzTLawBH74LgRpbFV5hVU8R7eLDXH/5nkJ0xy3Qv4QsU09VMfP37lEGe
9lGOQZ+fhuC9Y0grLk5JwBN1nIo+LlWzg6eBK16se7Liom+ZhrV2VZT8kEhzIwRHo5vcxmSmtYE1
N2BhsidcaXGWpy5iQimmN8JPGozqElC3dNYuaDx+E1bfb5r3VWte+9ZipULkqjewfpJOgYc95XyM
DRSiYZiUq3+Wgrhslwet80fdfYXGrwySjfWii7UMn7KFvgah7lLlcaratPTNHZPyQof4utyaHota
XE7ZPJjMT13yaS4+gy6yX+6tX7/4k6/TyM5tORPQoL/yYw+uIdSonbCGVPWDNl6LktBu0JLhIguU
O0gdiMC3K8F/1GPL9sSg0xJmU2ge6k9iygwou/PzOKXnHuPY1BMidCexb+/wG7Moon+GyS51vcfI
urxCfBh6TFgaI0Dp3eXNTBdYghDW6WyRt+sLSgJCcmSEN0+WmM/c7BnYMa1Wt37lzRHCRFrWHr04
28UXEa0x+D5PomCeZSxNRnxQaqQ0eO/Lm8CbTduvuvPQs7BCB/2EoDGRuGn58EBZ3zXhPhAvnZls
2te2UH16+7YCwPZCZaredADyrA/6xQppkirt04iWmgtByglAEHOgbAamyo9Jx3uriBgTV5vJsm9M
H3dHdadwNNlk6zkEMlz0WkKTK+hPL9Q5y8I4S0hiWVLh7dTN8g8BM5mWh3xw7ki1STjcobdcQp1K
RvRf2/LFph01OYaD8cat9s/hiYKBZNWDV2QqjsP/t8jCw8yT7LDQf38bppPhdexif+5XMzCZ88TB
w6Dp7N+MBWdQYC+4a6KEy7caQNEY2l1oJqXF7H2424nNTfNg5lj1moQFFWIt/g//UPWeiEjIgRgh
RZkhCBiBJcbL/x9dXtQ/m8UmelqUrxqFJWZMh4Pcda5UgMpVjMWcZwGmx/TVj1jRzGPSEIFm9B1k
Za2bvfcFYOE+qF8cTxzmK9zhPHJSMmqXpgX0gCDBLEevsNnzQ3IDRQnvPsRlvxQGFHl2YlhJb64w
/emkAKXka7/WcMilNIFeOU3/LFANm1AxRx/axJDkWj/9pg+xsuKOCT3Q3SOhA52faEjbBukU5nAh
PHHz9m2b6PG5HvNyejmPdbaXM1FK3s4CtjpKLI8kxZPM/y9cV96NUp/7+wcdZJgOgVUBnMjwaXC3
feECNx/GsFQf8+/QYnKGyoSZyBZENEty2Ibnv5vuvCiFMqqxdEY9bfHAiaRXu6kX1cck7f+kktpK
j8Lchv3iDM/ITdFkq7I4yJx3ZMw4oLLMZrq4aJmXw1Qu7J51Pe+zfkY0q6zv3l98anHEHqu2ge/6
286De2enevwGoS2zPBKKPWfomFFUFv/0gnHVX/Fznn9yO4oOV+hV2PBnxrddQ/wxSM5qznLzhdIA
qk1qOaEDy/si/7xfNI0f61tidTi+VyAbKuCDsjvhv9SzyJWYfhDHeSz1VFFF7BDyfcxOmrXkevSI
YEfHYkv0IhV8QEiYp69qokGKC5LBVvNPL1bwnoK5+oMy5Qp8zvPv45WIdtWPzqBwJqxXEzz2M/nO
uOuFUcHrGGQa8T4RNHLSSVHN3GLPstAIb7iS57fTATD98NsiSuhw9dcrP3vqFZli3JyxM7UjJoKC
UAILxhX3/s1mLemeMb+pt3WCeqqZRvRi7jP7T8gIGlyUo0rLMhrHYyUgItEb8q5PnPUopJZwXBUs
QdceI8U+qr96+DUIZSVLx8kNPD8ur5liZ8ZpExREfF9NPgXyaK/EX3rF3bFwc2IRptLpTzb07HM5
b/zzy2W4YEAsEdQxOBdXU139JxBiBbfN/L9c14A883RW5BjZnLu+/uiQSI6uLGvEScpdLY3SEE+b
ZIs7glDphyYKpT77IqmRxhS50Fp+mCWlPsqQX9zgXack53+77wxfHc7ywEVf8BNDHyGDpUgA4EW6
SqwKmh8Xwi0hna432pV4hLHCAemHG8ukPdZNI85TSkZke221opc43AOJM77ffYb91XKw+ij6QYtz
6eLnmgigcHyfKnUYyg7FDJmYu6aoQCM1cS1oMeFpIwf7OGstCZr6hQ3SH4xMDKVGQuQ97Q9T+H6v
FxSmRsqKhr+6F+mBVd167BgRI8IQUgcm3mmgUsZzs0RfmenL25b7ZbWgBKKrmxH7HGJDi8wtLtUX
pZytJcHU16awFEaImF4UNASSAQS0wmp1J+eHHfeI2rBMqANwUdK+mSKehLbCNAqzb6lJW41y4U0g
vRzXoY6kxkE85h2LWqPek5k17FFJUfTPE3qrz5+w+HMsofGmHBW0ey1+ZrVHAuaQjO3A4cpiZSqH
zl4BGmfIZM3SbKfO/qzw082mOXpMaJP/BKdJ6gmecjNomWPMP7ITBTOnPagbXwg/mFC5QfWNenJa
jdG9EfsAvFZb/2VzqKov7G//qbCNqySrAeJDeYIZE7clwEC19VVp2Pgn0F//GVkXI4LuMXyGuUaM
TsthIrX9yQy2ICsfn8xScYGGlRNN7PCkoeUcwwanAgNZ3xkv6XmCGJnOlVI6PjoR6mxVDt/NDen3
vN9dbPHWePB1pFC98tcOR4oAJHwAGi2qHrSFHmZIDxTCTy1k6pI7NSQaUogkKvEN8XGrF6naTeUe
yPMa7blKd2v14OOM/Adtm0+AtRm7JQ74gXVYdr+f5g2cr3jmgSJkT3l4d5flovvr4GLW3QuVdx2L
Du2+SErS+1zfiBzhzxqvbyPhy0FotmBZXjRFb13zBI1SRAcCMW5BPk+V87lNrBQiLCEVEqKKxdhG
nZu4I/DHdiJSGYUfg+5/eOlUT83qhm1/UUtYlbKKaoAv2yhCsDq6l/kpDLFhsM2b54+jWD9YyKT0
12kjJzrXEklnQdpWp4x1VM/PWz95dPHxIKv+bXQaM/GZfMBkSZ4xoQaoltz9L3pP2VCtXKuVw3oB
iqpwPWd9QU4CRw6AHOKLjK2qjZWyCCaYIFOAXxKIbbTWXBQyMtbCKqYz3aiZHNm6diejjPJtZBqi
EJk95iWFyBg4j15igrT1zyaW7VesPMgAG+xUWU0HgjAcQb6DnLDQ6vynzswxIMmEbpIIpxBuXAT5
yJDBJEfD60kcNmM6500K5jzJxh/iiMJ6ASMf5haV8xoRscHKfFYDIZDOmdxjaBXvgpzQzNqEim9q
qT/kMvrvHQy3wDQ8q2Kc26yDlacOdZ9qwtBNgTNAgpkpHhlhRkCzFLUnBvEs0VW8+WVxhS4sGlKR
Up9pr7d6cb7d503aTNJG05kzgUj2vfna8ZNnR193wS36ZhlMhrm5hBBFB2AvVbKJ7RrpRg3SEXLo
dzVFYU4Zw9Sg9RSdhHYDgzdBI41EHF3EsmWtlGxzRJ9tveTcKxON0e+O50jBbQVX2JRdYanMjNWv
fQXtwUbJUzyxubLIgrnoO7AIMvIPeg3AX1F1i69qlcWWSPKU9PialhCfWRaAFGXxL7A/7ZOOI+oT
Vt2hcD//0z5II/sAeqjYIbrMr8hQ7Xq9iETuGXFDlkLkLVdSp8W1EEB5vVHlzfTAtF2WI3Cyl9wH
r3jdHOeWCT20oqU98JPyWjS1oQF2LFLQqtUYy9TQmHd92YG2mU3IHIpRAFLp46wamxLD1Y7osFsY
vZQHQin/IpW9Inrwx0cylB09qpFQ1lnJSg7mq130gEk7rl6htNNQVSsYT8Qj9mGEeaZZ4gr6yjH/
P/gbVKybahtkfgnKMzOHvq+gawyUAkS7aUCYf9RyNECZs1xTz3tTqBmopBl+oUa4lrvOFt2ZQ1yH
pEqmd9Cm8DXKPchDIrezIx/v9/fnvw+ZOiguCeuqzb7kTNh4Xpm6C8pEFM0h+Xzz3T9mfqqHYqCR
fcV8JGk0M4X+/E2/v1vtOU1Fle2EqUsD+2ME9dN25kQhqoMzpVhICwrBa0571ufv+kH2vcE3TqB7
x0l2CCQSJNjgnT+H+TPDxX9AiUge++YrlLNKNOZyGPH+fVu9u6ary4o8ytv+lIu/TcZSktGi6BNw
xZwOEufup3erT004+W5+7xU1GsjLwYN22T+vQUnM1K5xLViaiCuB1xcwT44Ib5Ctv9yNS7kS9m3c
4PcgJ4MNKVL4NYOIx/wlRAoNRUYZvJgorOE3EHD0HXPA2deF1LldqruWYkxh2swa1SlbBDPy5tzr
10YXRjKRjHHS+Qjezbps4G3X1pXOcgSFyDOf/1Iuadnoiv0yuEzKNcuI4Ig1zKEGyMcXUq4ckFAl
kbpst6qGoljSiKmEPxU4vNeN428nZs2M3IUaV/ggsXmhZnEaMjngfaHLKg16PnwfAttB0+kcWDHb
yDC5HyHvBSCY1/9QocS9bh9JdHLNZziuwEfMfY2XJUFEqAomW28VFF0ywYicWMNfXeoCFLml05Bg
jgv2naBGYjtMZjVOO5KP+u4iispjVq1Y58vcB9m6RjV3N/zI+46vGRRyoPqrIQh2G2qvh5Hwh4Sz
OcM6Gwp7acPbP/QMN+BPUVjRrQFIzJoI+M9cbIZ6B7ZhNLDC1Amo+HHx6DJcPnTJNI1WXy2aVCpJ
mTXhTGaFFu8YTKdobOS2bW+mUYvmFyoEXC7Gzloy7YYDnuEG4NtReUigG8g30Q5/ZlNohqS/W8Fe
pH3oEcilrzJOUno6fDlJIuz+CAv0w7g6xnu/dYwxyNgacKPiBHImyNfdMmqW9InlI77ldBiK+Gzp
9FrMU0sPnqYi+ZD0pzM5e081//vPVIkxwXJQ6Y11X1L87CBgjOSj9iJ6wDePmVq2f0jKVOyl/aZJ
3rGXRlcxk1gQFZ1ydvT6WaqmQPLPRa/zjpZafTSCDlvYFpCHL7lnM1royxsDd8A3YbZe73HgNF1l
PYnFVFxy60atrOJMrPRZCaZXwxl54xIjk01YbMBvy6VfXV2TJSDvV5ld99shEuFmvjyA3oFUt2Jl
Z+UdJsSV70vj2I25YDgAAbNlIqEYiXzD6Rh18W4dwFbkxsJI+0a8m24RXhYT9iDta4J4Rqe7OVYY
DwtX2aMreRQNSwM9BYeJvcXdUDnHSBjsBHn87QwJYO8t+oZLRn+04H4VUYr4RbBdycGYJqJxcJZ3
JxR9GeQZTelHdvDe+Redn1nfg0gdgF601KV469nXUS+tIphX9WcxD+wXE2/6+fN5YVFRCl7cBB0H
YtFiXEcCeFPxgkri2iNFbPjGqCxE5lI+Rv8Zll+jLr3UKLN4dqhDOaVsH4SJvjDbPFI3TPIj/g96
MdvqcTT8g8smwz6/x5HJ93mUxDb/NokpXbhn6pcF0kIe9r3t7Hyz0I91Mu0bJUVqkPgQlo8RWJZJ
GQGgGhPG1wWKTB6/usCm3hw7tfbZfDz/YM3f74nODrLwS8Fk+mx3tXMPTDUcqAfpUMOtw9ILEEoU
RwBM4k3qh7Q8Aqaw1TuhhnJx7N6IkQ/Dpgjmhy1i+LK+RtGdBfd/v23te5G+kRj8S0vGNH/QG09t
PJMQ4rsaUeRySp+kDIZVC8zUVYiBIFuPswcgNmhpmy1j43XT5fgLDBm+FNVRwIRSi5lzFpySiNTj
Da3Yx5yY7gDkurm+fczu7DCkNlryV5WbWqzp2s4Y5yN0+4jWFJTFxOLTjydsOOADb9K3TiCDORoT
yIVLAuywNZgEYeYqbRY+UtcMfGbV21hGAMDkhY/oZtyLeqtRKnVDf7YOqaLJPdxSpXlwa2hH1hYs
M/dT0HA6jsV+6eEditx/xFI/yYl8+IcSow3hNFp9COkviQ/v5WjC9LQeeEkvJ4WEn8iumJxE3Vaz
W0PGH2mivvIuLcYzhZaVOpanxVAD5IvVtYfq2DZ/BFVvAWnoRbeaNSkI9X76+Ci2teY1Iie5CcYK
wLByA71zTB+nm4JLy2BBzn0jHff+8rl+p0OrRnoihS9S500JB1/NSKlYJlfkX4fA9Y2YMJTgR1AK
120bbWT7lyW5vla5ZqktdncmoNczVMYLjgghoU8y9bmOich+ZClv11aR9/mzmyE3rBacZONEAALD
HTfix8OpvGtmDje/9KJm/JB6XGkPFOWA1ON1NDOANB5AZV6X5Hk+2RFeaZ+xjdfa652o3MNyWMTa
7gkiUXKGT8cmoZ69Pn9Rn196PNvWV1UmUbfsJu5Z7/t4DYgeEQTmbeYUWzQ6BORrGnnuRb20ERn4
ALVj/gJsz5ti+LsUfeWKQLlGisH6FPOTP2mOZgWY/bl6x0NrTvID+0p+Qw5VXlrvFtG4KMOcpswR
GxSE9XiX5JoiRWIcRwJAIeIOQ5tL179MeGeEyDo6wGIlMeSKkh/j4Q2wEfHxTibJZDAd/TXsqydy
USjdw9vJBPKbcYTXg4Yzj83O0E8p+S+nPD+maVdYt4ENGvY2DhRv0WGmFq1ajK0UfrEFHq3L9EfP
PAgzCVubMyp9liGSH3fF2lf/K2sO3OWHHecKZ9judu5PlksU3fgpD+0WxCjsiCz9vMfFuB7giEyy
HEOOukQwPEyN2UtOBqdmIEDIaMHN5/qmF3A4k5CpODU2DBmLG2ilvTnUs+wrKN1VEDko/PG0u2NZ
IIpeXpyWhFJiA07V4F/xga9RIxoIpTbv7vLJQmptKD+8hAO0thKy9+G4o/AIAbTG1PxEBV7yfXvZ
74HzlUVkwQ/jTcPTXx7CgI94bqwGLbrMge6cGEqycA67WhZtS/tF8RLkJNnO4/GXgvfDEE+JWE0B
YOrTfqAyXswAS8VoIsN/fq5iXnBhe7EipwhRKmwo+qe/gjDAg/A3ZZ3TcAkeMI1+xf8Dk0q00Tgt
F/lPlDAswAzgAMxq79eZJxBu7+xLjwEyWQuwwlS5vQEjbmSkOSdcJO7mrVHg5plCXznGubQ1TFMg
qcIAd+3B5iJY9rHv+E4iAzUF+0XCXWKiTdFE3tl9fQ06ZZ7aNNeN/SP8PK96LBpI0h0uep7jqC1l
8yvHKwq9HeQtOazyP9stEHh2o2vdrIcv0AIGdU1+eA6rW2Yz8/x0lqKRg63Z+Uh9F//fNvWvmJUi
E0X65c+JDT4a57s90upwQv/kIVMewipGmhefTR2QBJgDd5BHIAe7x4t6LLkteOAIMqgRp5r7DgYI
WdWx3gx5/d4zgQtskJFh7Mj38gaYavMH2kjjAI4+MTeJbTE6/jG6ipsAQZk/s7hrbzJZT2BEgo7X
TnrHmPqXdzOXAyKh/6JdfjpA6xPLVTHyP0bw8h8aLrZlxf2bNZ7+jrctWbfyHlcThs2KamnO4cZj
oR33958ZK+ULDKU9rDhOhoh952Sqgc3a8Qcnoh3Q5Q/RW1Y367HhlwIErVbCYpAV+K/ybvn/gzp6
csiqj30JAbUGmDJCIdhSZmpG7DI/Z6FEcvvlsUtKnX78n5QquaQD4Urip9tJ8salf0uGSJst8flI
Yk9FvPQqRwEzDqrs2IRbcm3m2jjVFewvPG4CkThcLwYH7lCq48KeAjjCakWYck49bB9cqe22xiNe
4Si2x+nEAti5uYzdKBUsu76onLoPOYDFOpS4XhwVnKtQ68XRj/eZHXmWxb3s0rqiZvOfAXDjGhDK
4FLjmsUPi2mCGYKqfZiDy68rnOROF48kBo0FCc+wGxPlUXkfkj9a2wRh193RLraf8B1M3FChahYG
fGhilSe6n58KTQwDVC0Ns5RuunCwb9C2nns0jJEm8W1rShcurVBzSBy9zjO0QESQPbTxQEKcvOlT
DiGXChnNLD+CWzb2qjwURUX7wm4Kh1lDRdKSrf7FkzXOtF/7j9mIWrKmEsMbIb3qdD+D5p16zxo7
PPG+8D2MDUXLtUC+xdA/NT6Mvar09BPNC0v0ndEHD7QAQz2ie1x5yfVTCtVpLrU4sqjzdsmgLPkA
t+znQ346bO8/Bwar+dW5cahUNkONuyy2NVEUbJLjZogfIhN2tb8Ib6n/2UmPh7q+OSOuENaWLNyn
1FKCbllkhSai/+kVVj/fgRHMV9clbi6eKmh1PASTd+07JZFsc1k3Yk3i0hw8rlxb9VnrDZP96SfT
fnWSc8le+7QNyGJ1b9fz8JP8Ld9Qh1ORarXl4HiMOKH1RKlOPJQo0sYhVYgBd47eIgEj+W6JV73l
vg5PiFxo+74fpCD0jpZMiotkwri0rCw8T71ts3L9/w==
`protect end_protected
