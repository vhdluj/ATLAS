`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XYirKV07sZAfwzgaJMM4/Q/0RuK9B5xIhAzspuA2CLxku0ybcCqYEN4l4Sp08pAXEEGUm0mo8QDX
aoNF8VHjcw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i6AngR115DjQfCMLZqCPMygJS/hHKBNfRSuxEppDvG6GAjfB5MS9di5G6njMg5V5KCufBgOicmAy
+ZzznVlqB72PVhupl3QxL/LVkznaUU2AiCI+hmoQ1Qm7K6RukcyforW7Ct4LX/lH+JEEsclnlUiB
iJcQSnENiuQFRR5By2M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ah8VcQdLT7D3hmUmqZ/ymjuDSqAmpohOpAiFSNRmLoB4AOCTaB4yCTx/U4RsYmnMO1kVE59QRG88
jZaYl5Tooz7IfSF6uMrFg7QM148hWvD/+3wrrLGTzum5xmE50Rzv5NpTcXXuC6nKmFrqPJ26E4yw
Wp0wPC2a7DK/cSaEGRwfxTnRQY++DJkELvDGbOwfEUYs1JxVusx6Tjg5qD8kaIAxoR6duacgmvTS
rythzOwMJIco98Fbz8ctzizahsSMRyJ4AJua22pGIFo2xIydKhdYqiQvs8trjgV2lOJAvbSyGgrY
HUmW4CzD7Ccyk+p0hwxVUtLLnI3XmF2ANJQ51g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3NYKHa+IfAl0ZlL6anCxfHoF9nungFuaPgfOUtK2ThADh0NH8zxs89dqrlDwT2MfHYI73ZOTfgQz
q3UhpKxYFBQ5qiydMmzaBtBL0d8rmVD2hj3APHkRnZnaK18Xwg+/08k7JW/GBJBXQfGnx2DIMUtf
1Muz1zGF9O8rxyOiuoc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FjFR0RvsZHQX9Av2r4N/A7PQKTjDpkyOyfOBBLohibtW+rO1zhnoRd010R6i6ndlAiEbl6xmZY2D
Vspzpb/R7FHpNK7MDYgBCmkzVbeVOg4jBBDG9WAhA7V7iqqRpkHOAkOzM4WjjK+LxelqqZqFmcCl
c4bR+bxUrrjAYmFQsU9+z1YbSS5ce7GIfJdmuDk63+YMsxMqlSHjv+Vtmoc7WeiUWmGYWWS7fY9g
sHl6XZsjLwEyPjx70GpfKbT37jCDrD6Zxz1/Od2RF4KXhI/gG69JegfaVawSb5zxU3KI4ZLUlV4E
meFvdWq//TP2F60qDQA1fnPUMgQJFsQbY0tWeQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28400)
`protect data_block
OZukfODx/rdpZJOORTyH5rjXKpBORhc3vRJujHfOU/oebL+Dp1TALIIsK/8tncl5GFMReSPUTcTf
FCs2KQ1G0eQmSVSUb+C6jZFUTLgFpQWMEnvx8Ki8k0W4YBBNqkUE/EAg3zdEgn3YYwD1mKvb7o/G
yvbK62k8iBXhvRLsiQvrm4m7VgxIHldob9Rm0KOe8+lp1SbJFI4KEYLoZ0cMNzMkGwF5WNaPveD0
twuRePgsbaFfkBUvXu6rDUQLNUoeisi6RHmFicbXmRInxrXX3Ur4W6K7atz6tcpBP+CxBYID6+81
GsKEcQx4PM7bB3mJts/6nH05i1MAkiK01or9xoWs+8irEbvxC/28BnJeejueWOfl/nTTTcmxKMSA
ls71DHZx6n0YMDtIJozmlJmvpMmU5AkJQJSJf1xRSc3wySqd+rC2Ey5R1QmcY8gh50dPTlsX/YF+
C/D8h895tpuXGSiwTT91uf0VfBH8mkpEz52HetOYI4c94PCA9wE9BR3osJo1Sm7eB5ZjP9A10ljF
KcaoEWzEoafsv2hx8FcDrxUdT2mMnMLoWhpoaQWgGE5MFZzzbEC6waqpntLCGKcpwDHv4CD5cwWF
nDCLT9C4g26HllA3mjV7NGl/JM0p/SZKN8OVixv52j41PPFzKOB585gp9CP31wIUCFFY746PkMfs
kpY3/8pwsJ8Rm+zqh7wgS1NHwEPraPAe99P4ItaNiILgZ29L3LOabP3jbkxm0pqTb9jsvoK5ahs0
WpNBmiCb/mWdS7TD6RVD6tJ1uTIf03yQ+jnSRFtqa1tJ8PqcSYWdFi+BVciG8ZX4u7pgEzf+j3cV
F1fvqL8vwGv8bziTxqW6jxJi+QmGPdYR4gBHgN0wC7IM+rxCm1Uy6buT/A82zKcJmQSZEV+BNzFt
ihDDbWngLrL7wWoZzpUPYFXobj05tAbVV6doLS0mkm4988mLYNJvPFWdbHI6W0vV5j3hEjmE6ywu
I05KbqFMCV71M//JUdDOHY/9lwDbvszQDvdAbas7QonKkFt1wDWh2e9PERJtms8URqwk8DUpHZMF
0B2icI9SDqCHllZg9+IfGkSz/zF2iuIYchRKA3TDLu2K3S7pBFDO0wMlJ0J8qzNSFYRr5DJdMBc4
8c+/jWzp7X9BrdCc2ULa71HQkoosB949FwtSWhVnGPJiZCx8IgKJ5aSrLFuCweH8nHUR9Jo5BSX4
u1qU3Dl+q+PNGFFsA7Essyr2CWy7wfredJFEURRNIElIK4K4DZbP3BfS06YMgJpLXUj7XwKfbw1U
948fC+h6nYALehcfCbKcQaB0XrIcfVpvjoeQ2wkPsCCHsXTIm+n/T8A66lh5RWOV48iaFhJ9mt8V
8LnjcpouQIwu6aeQi9TAPdFIfXi4LLTuRjASAaGIeky5W2g61aMBiWZJeJaEeSQWB4JzKghLg696
cBsKpHhEnipO0J6V3ivvI53NmJvoontfdHAFi5+JSQKx0ak2qgJrZkauz831wcBVl8vF2s1vRT6R
/lUJ+jx7BmbvGiUPLOa4BOaQVStPeXLSVFaRtKqYxc8IHWGbEXbotqvNZTygTtirWi8+TH2tgCxw
MctVfNCfb2LiDEib0y4OlsKOgtrs6bDPdYn7W0Q8TLauivxeYImOrrIoNR6OgfIqLVnejt1XKZz0
KFgt+6Pt0C619BBDAHCc+jpYE7VLUVcoFPWJkpkfQNDHRlcqefISCrSMaeSPeB62GBdhJ4yW7QWp
wjSNN3PmeQCivTi/E/zy+U33u4GodoQR9/G4JMS4HBTsBV7WOR2VoEI4TaDEmXeUNdfp3ODlDypF
GC8nUqhlzWh6Xw6BLFWleAe4dzGRW3wIV/cb+A78bNXieDzuQqaZXcl75BL9WtOMBv+nsyelzT4O
V4qUSURqfHPtqZMrWziOdVuBpoU7t4w48o418ctzSR8c+IC8asSoueH+ubN0Ww/ssM3ZEwcAlhPW
ptUjz0CeAM7FUf++VUpyRZ5BMc3kI25OT+RckmSYdDjCtB9uolUMolPqBdsgxjoBXqw7AQWFGSph
XmARXZyucCFNFhA9tgiraKLecBVyQcqZ46t0GcKYduHWvJb/q+0V0UxdI4IAiF97aGif0uF+WeCZ
DYQM0z7fFnAd+7aNvl/Di2Lvlr+CaCsmXradLZiCiNWIp2oKWnpZqVSHzsPxlvB/bsqFORkCF8xq
PX12i1/GptHXaP21g7rnRJKZ+tvnrsKT5Sg6oAOPajkowtWShohiSm1Wfo4cCHWJKx06ngWDhxON
bneMB+iTn094iWRdQhehdT0l5Wm0BgmzbDexLZr2omWsaAaZVGKtMiLbwDtMzHM2kQmTlQiKSRKP
IWvvRP2Rl6BSNAP/29xnT16dTPu3NRtJA4K/vcWX37WMtj0hyxD1gbq6s1rzqKIo7rz+RB87naWm
XT0wMz+nw/ZTlL2K9xrcrAz5yas9Or4MLH0YhUKt8UEQX6NAWiRL73skiJ5Vl6zHHCjgYVda2n89
IGqHXcmQkZf08wNRl8XxToutI7oskskOj1uGZCpM5cW6ulkGkZz77wwBoMmE0ei5Y7GYXhj3QdhC
x/xHHmtg3cietrgExxqkcQG4V3b9mdxzpv57LWosrwb6mQslaxz0EKqZ5p0voq+fWrhQRbTuzsbp
ElDegbE3FDmpTCSk5iup6rigcmsZN8H9Xl+L7DuUbmUZEQwVjiFsU8Raf3njO//RH+fuoLbGZD8Y
i53P7uxvmHkdiQrXoudn8ROXj064zwkeAqRkTNY0qhk62rrdjRp/e02QCYRrpOI0ZCuT0XPUPcR8
mBmT323qOU+946vxtbd1suI6xA/OkCO36Pc5kjU1h0XiVRsGgaR+JQO+x9b2sCAPotr827W92AYf
HPCfgoN94LCMNxHkySu2wRboEXPpzov5y/WDIqDkKdmGbI5gLTSfqhKgI3nwjWbjpgrlcO7pFAM3
6tWr4tAomxjekfMhE6ZymjFgF3ehLQC48Agf2GmZMBMEEMhZhtrTWgH4MezNpQq8/kmddmNVpgRS
SwNMfQDykAtuxoJx6mnGrqhpGceP8dqBqAUwNOrD0TyEfBapPBvlMDrchdHRWPE14f/tKhZrHOCn
tkklliKhDreD8rNwb4y2cJRcrWcSDZH3ifhsv7Fk4BddU2GSBBMEbjqlbsklB5EwHNKF6e7ejtYQ
jPhS5JNu6nCCFz6BvSTahe3rvqscm50EWNURoqDSjauZwkRVJOMOp3D1EAzHaN+VMujx3O4+DcG2
ryVk3IJh+0ZvYSG49b14Um7vmHsIL+vX81YVMTIGwvhYdbHeWHmZMrhXv6ePnKuOXi2tgVOrbizr
5F98QZB1MkRMAE5mcU2sh2VxJnX1hG1NIyoYHkyuhwAIEzsTJ9RYY8842SjilAinsUnXASudkxPz
ihcReo9y+wG5G/1KMK7zrEd7oFIfTE5qjdEGIvcZUjegf0h7uO+IJBl0qeiCcrvO+bNsSxkZaAUs
SSdfTb2g0V4GyHKd9C+UV5uVdyBCKQ0z2hTIacGWGrWZ4899O6aa2JdhRUmJ9vMjTivPKBsnpDxY
pR8JVh19pgo9qMP88ftx+g1y4tLTdWL89cuG6wuZFCpVDYzcm3k1x2JHZ5fwVDDQ4CGi2IFpOGbs
qged1Nj7O10zUmOJm/Hqa/Txe11nHbHgc27ZiF05iDiHwvf0/AZsSNVk/Fu4t08xWLsDViYYugxD
EfW0N33I6WTie8TdmKK8QrZ5qUgsBHf8GSHW0l3Pq31zo/xlgh0iVIjAUKX/l9KwMgYDlYiosU87
CBxHR5v0drtUK90d1w//6hOauaug0rHXOUPpFN8td5+G1DjoMTs66CElNS1tuP78as+eYhi6PZGl
Q7WBEDvoJ3SWdfvlTKz11UwJGYjdAzphH2Odv25Goql3CKaYyF3pK4AlXATJ2znotqDv0VyqMK1/
ha0AjC7BZSYu7NCe/xOxARMft3LCK8j3yDqVjZuE8O/DC//qZJ7zlV7IWeMuR+VCULuQMnGeBq6T
K/D93mn85w0a9nM7AwiHGvYBa5W91rlHerxSiFdetVNKXu5tuTOI0+0snlKALyU2vBcGhmcKUaJc
qIOOy3cex7UCOkCrKcV7jUn4dIfKedL6So78UcV7/ylVSjhNznvIub1PdQOOeGNYKJwf9i3t/4Ey
WJSWVwHhsadTRWpHP3Czz5XBWOFyvQ9ToVkwTMwBco/ywKwFFPsQJEOtCE5XQP7hf9KsoiJ2Aq9L
jPi8GrYQjaPMbyx+IWD571CQrE9BKEG/uk09XmwunD7Qc835k2Ad2h8UVhy5KlHbwe1zW6cWZVvy
Xqr9WYA33DL8XRjU/13+bihUMjP0XKLqIkv/nyjckMVc+ihT486GdeC7SvoSoNtQRdRZ3fQxkyvJ
HsU8CAN4lMlMUBJvPOQog1itDtSC/MP43no2Vp9CZYnTHtG4fluiyBE2ZCzU7ZrZLL33jTr17lof
XtBXG35S0S9PI7V1GmPVVUc2V6MfAj8+Eij5gDQvHnxWpbhpZbAIHdWw0I+KNa7Kxc95PccXXCV4
MpjHI5+lLFLLSzoCzpR5ve0VbKWY2TMJHo3p3N9b61J4Ztym7b+ushESZwh1sumk3QmC3HQqEzn9
j9l5gY1+CpOWoBc5ZKzHSd+pgww9C3wfZcKcehbgI3KL2iclMf5Oh6fu+wd3xB9U6qUbbSL8mV1o
Cyw6nDTblS2uoAK06qoWwl6bZ29tEmzVVXwAyxlxUJfuErAGScaENy4fdVT10Rc9pVQe2n825FlV
1AvZ0dXFGgFWNMDYG4BGEbQ53FWEr0o68LwRkVCkNrhlbF04+XjKQvoVhmHCqpYI8mz7tXFid/Pp
7z7Ph3WQY0w5ANrqS4REEeRNwWujvShEu/jij32fMSWv2i9Pq0KW0DAmwpE2GuWsREUNgBphQckD
sqAWPAcLEOXfpnU2K7x819iMnBTayvI/FztTWQtnMSDz2j1RggEnnLpJVKmRJ8zjJbcNh6tUZXa6
8WGog+wZGgXggR0YN6+SaQzHdEuF7TK7W55xfKLEhaC9iig6wbEH3TKY7TWnBfB+XLt1W7MjJOU7
SrMJ1Si6bp88FfN6H/fT/EEU9PJbwg3dL7eOIxVDPieYgeOC024vCsGLr3ZbJ7Oasn3oRTHayIL/
hjrF1uowqIEcYmunjsD+mOZ0mxS+m8Oem9JfhCGNG+nsuy0eTCD+765+bOKT4UT8oKhsIqvArI1Y
oE6Ltdxr0gIMDl4a/gffeEhPZ49Kw+2+SBMHFbOQeuVZx1cWlFmeeDhE4Fqn9dDKr3p4aX6SSP2q
QmcpVUcLnQK4fZvnmt/uqebue9cIk2C8PVwaU9M4KbhePcniwNrDtyzsrsGFoB9m5ePhQBKZ1Oq9
CyTSa0PFGIaquub78ETGXnPPnfUlcbAo8ARtl6ifs3DEUko+c23kaIup/d7gAz3evLaalPZbijhJ
NrJb/NR8hdJejhfXTh/gM0j9BBzhsClq5Olbq6QFb6nP7GzU9XHUtjF+2vK/u0DjDtSAiohJalog
ZfljkDIWvGxQOPoHwhsDCHF0j51zZ4M+7/b/25RAokkgb0cBHsEGkZVR4Yw4HYOZPa8FhZS16eDc
mC+KB2c9dEffX3FsSW/p+hGIvNUtTi97x5MdYn7nSUIxxjtKIs5Y3yd7OUYs+8UE3JpeMz4c3d58
PKpfJTct26sTZmjVXuU523kh2z5PAP/F5MiG85X/Af6yDhjMcep4krNBY30dFnwwbT1iG+KlJoIu
Ab3xcPgT9z/XegM7HaYXswS3P6/kSZqU1x2XJfqp7+X0gRghXsPYRC5TDxlwigbY2cKEXKJMBRL1
f1m7/GDVH8lsKPjzA5Ex7yV3OmGURijV20vJVOxwpL+84RlczWp2KWAS2dJZxngHDgK7KGO9ZAGV
VoUedRMQALLMnNHQL9x/aM4wwc99eoUeG5WUZjgVMd78wHZJkpCLzUxEK/OZObFKnJjZnae2+8IB
yCMti0ejQwuqwYcnQ25wD7XJtEVFGs3Pm1dVrrKMp4pTSUMYGMCLYXTsHS1H9AXyA2WhrqCoJ6q4
NpeE1T/RRqJlSMR5uFzYsxOIZ/REqfZ5bvHdezJyuqFH4FIBCluRcMBPWDVzY3McjvPVwySWmEJD
MdLbeXYfhIDPbYIJS4xxJiYtCYp3qZXgj/SEufYyrN3oaGjrL0mvJ+63uV40991SEZPWgXIyV2tu
+3CilD89qhqZ15KCV8iBjh/pmy/QIf95WuCZEEE82Ptw6+8P+r3k19LQp6pjBlJQ4mUJDpEE1IpR
gjFPDTd0VY/fvJv3fhJZ1ny6hClDE18RZZepXuVXBH51w9XYiwIDgy/+ljQZ8w7nbPD5E/dupefL
4G9BJ5rdpb3oNGpQFuyFXmx6uhURWiEVBNC+9kxacogp2JC+Qu1yCNIMraNKU2m6shtbAdqQ1uHe
xMj5Yzevtnzu8ezydtK60qs2TVRYUVTSajcT8bjrFhLqvhQPTMYIygHWSwc0Fq5l4gKVt7hlFzpP
q9t57mKK6Q78kiRsxT3P2rqwuc8Y0H8wC+iF5RL3xs6A/5GCd1tzczSAMFIY3hYb+gmjHBuzrc4G
iQ5gv4a8Tp+aQJ5cNkIxpwprhFOVEvjyYx2BFchWL+/HAPh5cElGfQLdJ81S7Wbnh3PM1NPyvLin
iIwSNGv+ze8bxF++oUx4MWeCxt6TYoS5YPF+Leyoy71PWcLLLQ7MRhiAgaAr1Hg3OWk/Q2tYiJ5F
nCIQckrOxV5WrVI3PHOEdgheWwgukR2f5LjYFPLM0j7835R9yia61qwJSVA93e1cUyr8tsbHr1/r
uuewYImEpaf34TPjy1SMtzy8iGjnpN/ryXz6ksfkD9v0XXNmIGnaFoaeQMRr+dPG4W0iswigbAQm
4pMTZjxBMo7o9XSgxAG13lC1btVIgA5gVDQqfV1IIk4m6iou5H3yjdmr4qG0U6yGMjKtwwnZCSwI
9Lfd233z/YbmS+G5XroI/unhR8aoPSzIVLgYC+fYW3HdDFQxuhTjpclXL2imHAziHu4ib08gBlxs
aY3IhzQ3azyXggw6cqMTiDnvpvcoW2YsmZIUHNJlUrdqRlxvOSH6/I1TiymIrXnesC3JmWtbMuPP
AiUFuQaXcyvyj1YrfKhdht099aV6qkwOHwYnXbrtqnXdOKg30TXR5Y7upWbRrcxFcLZifvy80fOq
8TVr1Knaw3FLgR8duDPg2KbrhVgZ7UuHStLWctc8pelPnuaiudl+P/RspcU2g+kNdO8juSOj+IIi
YlW9pTpuY/Ag9ZYhfxaafN3FT6M0Hr/1jyOnpibjjYuRcTE1PrXHve0Jqjq+5wmoKhOtGOtayeHA
cTZazDPEu1/F33KgWvKqVnn1852Y8GmbTcuah0Y5AHdoHBNLZE7sJoYCczwFZVRCEvCmTLP6neVv
GZTcJpgPcR8VYGEjWpkiWvtkQh/tYYN4sE/I++Y8BO1+gEjZJCodFFNWMIWraDB5SUXlRXV9598U
ilfpTe5nIWzn1ABe2KG+6nSCs8lwizARmj0XSWSSrZjtBkFvjpRUYeaZj/SO5OJCYE5duP43q/xK
j1xTxQZ61DRtPSfUC5Er4+Y7dQzMednYf8YZcsu99RMCP/eVhemyVXVKyiEkVWsXhkU8tsMcU2jr
GMob/cuut9GRzV1fwnmepQQJU6RGB/ziPXH6wzEgiOwjpZWniLmH1DgAICbu9EJTugb7bcdTjC22
wlwwmnlyqI6AFzRDtDYeFhF17meE0Qt3MsiRNnWPHwlRJHu69cnB41I3ExHWF7IT+MGtW/XIg76U
2FuDmiBAxGqQjCH+gm3zH0dk+XIQSyfh1kHGhzJohjUG1/pPPjXheb5Q++u3HE5Tvhh4y3RmHPXS
FhHh2WdGZHBZIiBxCVtW+ssLtj/T6o6Iy7AwXu4/xlyUFs1Ob9yl4uvLcFPyU/dAbIQOues3OPuJ
4pd0xpYlvI+ZXcYcOqvUL9BbkgrhgJ5Q/MVCxgmPcgplBTRHdfcuA7SbVcX+5N6oAOGoA9tnvYFR
Qi5vO7JHj9aMuLkKevGlgSAES5BfIv91Z/2B0SxRN2Cab0U2N0KpDEPJiL/bP/Zzcq/l1ew1CjUy
kifmMWM5VuXvFvHIckZDwjD+FGtZvYt+Lh13XUSjx0XSgpHA/9jdkoNcLCqVpZo13RY4yZfWNkW5
Akl2swgPqwKTVYiq6tVpvT0wUIHcFFhR/m4H8rAi6k87NmCMwWwCmSMjxHbQfwy5cdYtncJVY9dS
BIjzH9I2I4FGPXJCBzQ7PvfUE6jIXGM5pCERgU3qRZPItIi5ATSx/FI3xWzpr9fhywSYYlp0K30M
jknnq1fksYnOYK7LiBmHnn36GRKL2h9p8fqaRaHAoqMxBm16IE/LY6dyrkiOZ44iTels4r17sRgG
BIFGnp0Vrtm3vtg9+yIp7L7Vj1VGTyvR7Qpp3kKzyP98+oPZ9H07W2HbM4SSw9lzerFqUxhrSRMp
OELF64KyjyiAx/kfirYbf3q9yAAUjo4zxuFx2te2SE8spX+6e+a1I1I4oQuEUohxPxYg0tX8JAPB
RI/WTzCE7g3Wi0LD/tVJYS0NGbI8NpM4CEAPDNjF3TqNqemba6tQWhGG5kYqaDyTNTyqJBjBam5y
/aeBCXFZu1g2kxSyFWOre6dPJg3XNMIGE6QQwbxGKFkpv3GRQV42kBmj236IZ/ZdUKj0EtjChHpc
SguinrHs9e9RBLhhmFDjN+FE9jpBTvsjmj8KA7duRPfpYzHXhqwsrpc7S/iPxk/ksS6I4AdsYZR8
BUeWYZntLBuY4C/xmmJPnQqYzl0Fna9sY4ngr02JWCEKmdERvsOWGLKR10NA5AhHqYqjSgMOG+cF
VYJcxep9UrAdQ3/TvjY/lrktKTpeQP9iRrf9K9fW9bAWlZ6v+AQwuWaE39JWIxoftDU7DkPeeY58
dvkRV/+kKJ37iHEstqB9N1PkpV2IINaX5uP0FvQjAu4ujh70ahpA0hlyEjVEwxqwxWIan+zaSeZh
iwuEKvOpkOMrcoHoFlxO10isZX4jZ1DJZ2oMryRua3jtEXQxpRBlURa4bNvJkF2yk/IICUkJtBkg
VyU3RjycLqYzvUuFDUy5A1kAqdrH1Ou8wqCs1nNJ7E9I/ixAWbc0SpbSZW8UL+MdpN5dsQ1tP0kq
0XkliRcnpAmSFLAHI1Y5POGhcpYf1NZ9LjmlsLMwSYwrmfvnY5lSmLoZDmnycj/yMn9sm7GDnsOX
aJUuj+UuEOBKWcbIoziXJncRnTS8SgiePxPApUph8nxXX+KUzjWmaKIYlhPpHafB6sqUl1LKR1+c
4dBMFo8GtB7fJolhIpfh9LE3Q9rQmiB4W/HaN7y7S4I0b8fZI2HO6CYEQQs7h7QHXSotnUp5L9MZ
pdCtBkltwhfC2+dY357n7VwZoMEUV55fyQpVHm9qWQRXbIumsckkCF6yQNOyJvOkYYejIX1v+dVn
dypy3S+KiW23jb9IgyNGtSeZphnNwnlN/o+opuixFfPtsr+gjo81pO5LnyyvBeZdOJGr9gfUeXkL
7TdB6aUFIVndG/BXLsfdZdPTFq5qjU4YXkrFyIuh3hN0LX1MSzi/bVmIKQJn3UmvmMDwWGIrpeY5
Fp+f7mloIvHeYCNvKYwbOqpIl+rbB2h18TIf+rPAfhLuyQzXLCDO+osdrtR8PmRqAsYydfLT/vAE
vDE9Il2MCVtCBVzYrSERC5LqRFNSKlg9HPSDjEzvfEdpabHJcd8ueLTSDBwN5M4ir75nFhPXL/9u
Nsef7DjS5ZBLqBJr3hGtrnA0WfCkyHG8qPJuapgPGK4kUMi3ZZzMvjQlQAqz1gP2jALuUR2a/+zl
pvJbTj2UHbPWlLBVUTu3PbWF1FVT0C1OJoNiYnzCvV58gcR9sbMYsXCBkpH5xBTQzdchSQdOJBiG
4pZ5mKH5Z9LiVy13QNe3CUDw1GQ7GUPcj/04RZzhmWLfwy7I2OBLHxPf0x92FjRaBPBHicwUsMTk
1/fqaWQ/tLuYu9rmgy7NgttStXm/q/XWGPD5+w63DrdzKxquqVboRR9iCgqWdFah7sIFhVxJts8c
ZC0+28Kw351Ah4TD8fTtYyAoG6dFHn3JQ0f+YQ23IkVvzmZrkk1HTR1F5vz/TXFF8Qmtfd0e3GA1
auEQWEQDe432W5D0Tj/bDrLgIyCS6oKGLJAKJWgXEYAARWbwl5qqcnPDcYuYuN5fj04Nhkhngr2J
yEkW787ZpWtOzsKPRkFwxw6RSlRTF0esEczLOHeFfg8OwK8o2kepkxBLGOzxWJbPzlIbzyXI6R2H
TTZTfZ+/2A+6JRhV3Et2/BiAUPI0VNX0m9EdqXf5h87ZXwCFxuz9ccVPZsjuSKw2d2SK3FxfCK5R
N3Xp8k33GlUV6oFwUQZwTwnHx+DK5OpQIYaKLMB99kNowKQtEH6klir01p9eWhiVPexLC3edaOUS
7GfcMQ5rlCXhHp6SejBWXSRZjZkMCUeMAzpyCUSiZNVqs+TJokKtGjoebtqqOzZDU6nXcgnH3Tzn
+EGlwP1JK3b5Xlv40d9rzTfe3Upe8E+fyAgTN2ZceF/HbVq5jxtw4OmpG09MWNMLWT0PwLvQZjzj
f3OyFf0nDY98fYLKM4fXsZBa/esrWOhlgSot929UAFDdVwamatRLOXzlsypkrwWMH/iFbUxb1Q/8
B0zQ38uhvuwiWN6ApXhl7tXhvNKQDoJzbgM/kwWnq3yABcupZYG9xWvDijaUq2ZVhWQ9zBDtmolN
SokyXdDXRpJUAPPrFU2KEb2FhlAo5i7dvbnx89SlBl+iZRKEQEj7N6vaXUMUvgntZZovneWKxCIA
bcvKogeBHr9pAE5aAeEuhmlAByEef3zEWHdlMxNxzS8LlseJ66wtXHRZ9QnK1fSkxx04mb8zG5TS
TiN27U8NchlOEQ3FA7TMj6vl3fQv6x3ZZpVRdDj0PaGvon4KjEV/YIHgGcuCpMNSTCOpNUJ5teDR
fbOhyQuaHzN8KldrjgEONxxyCiaeSStNp2bTn09+eVLs1+P92Lp941Fgpa5zFggK6yNhPK5dG8sO
xabePOWfGULuVAFSWYFzNY6DMfmrVc5Z+qpTFdVLlvfdVpoY8JgPL22B2p7sFmbtkJIjB2biMlfg
ZUWcLEf7hZFwUggLaJCmRr9OiIL1lVlAoviuT2OqVv8st/Tx5XYNuAdgoDjToJpw6w9qvsZIlE1h
Tom+cnPFQsoIlNvirLfsTpmcRuafxuNVXtzXCSZZcHG+2YNIg4YH+lAQbHe/8f/aEHVPJ7t3PiAu
hDPYnB/ShgkpAyCrppZgVgEGFO98ZhBIrQ8SqcQVb5pnpnuBUkcoTUE0VNCVN4cisNKIiQLUzO6A
gq6LzC4PCuH37CF5gkH8ZPhTBBWf4yhs7YDhetoWIS0ATFjsg4nQs235EeVdMSBMuexBlycxAeh+
a8cIaGC/rhrTNgxFAbTGecxCgYTBplKDjZUhQxnXeXwX1h/I8JgbncfpGWsnto6bCh4IfZX6Oa9U
AO/rUBWvG94jiSu9sYmR9T0p8Z53e84oV4zo/mLa1a6bs80b7KcrIQDpGTV8Y70Y+t68sZZavdev
/cB2Afy9qMNaCRSNJ+r49kaD/iFkXjEtPEQxTr92Z/JbkaiHn/Co9+oal/UiB6NuInf/Kp7WxvZo
uv3G8pDhHBTHqxoayOgAr0o+filMe8LbGO9stuyysYUUA2tVPBIhNWdWvl+rZrEQndjWErXbIarQ
95EcZ5taL3y2K0Y99F7Vbv4zb42qCRCd0hnHQnHykGKoHSa3VdwY/bKjMl4jN9ICBGfNxNOYRznE
7a74k3+2y7/KQG7DdK+XfJz27YrCMbCH4JZu5rprcahWnp6C8JRTzBIQlJcOQtkGWXfGTXK70b5j
saJrJ9yVaIXAgMQCmWLLx0u2/rSCt5EGsmfYkx2cMRl1jJHLAGGXV9z9Ux2ttJg9ZXqXnJ2oElpq
o+Ypl2Mnq2qVweQms3RjltmlB8Rk/Szix6WAqXDvVHa6JpxgCH3vlO+jyVIu7D+MBuTFa6llp+mC
YgL8PF7C+lhUdR9HXNoqxak4Klvc7wZjQyGjMH4kfnaSN9H/A6ysntiDPWuRibhWhT4qIuSlrTwe
5AefjFUfO0o/TrJSmO47oBoYzS5lkMH0T/tsB0FS9yFpEYYlfWrVBS6e1yWnRxDva9SWQm8D0LHu
x6+WFV73LutD1hH9UIUmSnM5Ibb/fc2lQqkjh+fDbsmEosaz4Q6zMCyOzdRiztFwQoFujoaj4KTB
8yZbzn94e8FsuJWiQ/r4OelJt+eVs+/kXxEYV0O9U8Gx43vttTAaY+X9HuTH5DhYoKjlnQxHw2Fk
aQElAO03A6ZwpA8sAjAfqjcDCrhazAQ9vTY93dEfClm68LQIu1J7siY21xfqE61ZrBnWBtTWNadn
LRdvGWkaJGrF1BQTCh8S2LrWknu5kfTw6sLNX2rJBzCKkfwxoW4wZDWhc18hEe4aRdylwVEhHrJn
kqrNTRFA/KWZaboh+0mbsu7hkzC1/BounfHQRVQ/6JkbTlBKhb/AbaKyGpABUbR5PrAz0cl+fis9
hoc23U9w0aphsAt9leqetq0lpTMdfTRT9GPUYgXpe0JJrbOuQZaL3xcpUyZemSiC36xc8P3wWKrV
K/D0NlziW7t3kUV/fduE8x8fdDdNQCQIPEZsZZ+TfUeO7UaaAFzPTemtHupR7JKeMtN6W/Fd/ErB
7+O0FNbJHU3iFqX7Q/aKre9r+NNWJQDWuU3Cpu+XZeuk9Sk9C0pXdzFFp4GDi8azq3JIoNPX2//w
cT2uaJwL4IWYBaak1ZwlNRBdRmI7J2SGwOzli7+7iGrxC7b0oja7hva6BYD/DWLzgualqFxJXv5M
YyONwxp61Fh2GpKQavo7tru7fMtQxvDJZM7IIfuzNnj6AK8YF31N0jY87w6eMtn4KNHq6fhnm7y6
jm8Hk11c0w2r4ASeJxq2xkL/6rn1sgWmZBsyro2lsGzvAQ8hJNDrGEX4yADyk5TKfPFAYXWJcWNc
iBQB2FdhEfBkjlku9Qqm9PGtwT340BXETRA6f55ijiY+hdzvmShD3+qgL1jw8woNuJU3R1WuN7hw
2Vut9bDgIHe630GsRYnmENqbu6+zGtiRmdxub8P+Wo4UxJXR8XkIGC+ft0wA6UpPq0q56tYDKqi2
7pgLCR1sjvODg8pH3nnJ16VaVpvvNj9JhZYaL2b61wsbbWV9x4rSwycmgR8fWeonfGXtoQKEAOkC
fEH7/BhuZPgHar79y6FnhxuCcwiG+BaV27lbMTaJk/QLJGcc7p429E6R23Ke8oqVwge0QCW7qGEh
G4seXSlXpS/eCEGXT6yls1VWxFgCoUxPsQvek+F11HfI+KoVVM9L5bKv+5dVt1UWjDyhTdNa5HVJ
xMBkoQCtmRPZ/ZaEmKLK7XN5PMyAJqSii6/ULcV2WtOmWRneAN0thU3KWjBJ5+PL+Fs15sC92OdK
AeiLbhi0qRIq2vOhEWzZpz+sJZ2b9RuXfZc33cOZf9R5aL/XLrYF1nnJF+YZkW1bxm6fvqDodifl
2fu/OdThRmjOiBf0cZkgSfKlMxYfXua0at7jFMIWR6rkQ0xhAwmAIJfqSYjfWJn/LVN55SgkGH+c
uaw/4o5Z51WoMYyzN6d+8jRetkmKANLadGAsqRGLMWvANaB1tR8xR/gFouyOSparAfdumYQsdcce
nabHYtAe/yJXs+kiAtXW7pzr5mCW9ZB2YVyNf95C784Bpxwc0x/sH9I627G9KRYzrzUZ87EHn/wz
kip+v8mEeXpwolUP+g8MDpSxlvtpXqCd3oARRH7SgtH0naVxdIeQXc92nddl0dDWd95pzaDpwkE8
NPMI4HzRgd1lTTBT3zVmr1Djv3Rt2N8W0Vr2kZkc1qwU7ye9MbK8s99UPKi2J/GlCorbvIY0R6X2
F7Ha0sdnQ2GgiOEfWgB3ZDYBG52bJZj2OPCOCqxMMoMfEfUUsIRl95303S2yll8WkCdmiunYYIZR
ll3h5rH2gWuJNjlId7+Kgh341q7jtRACCOcVSYa0YJCLNS+jxUlR8qGNivHHLPKB4+Fklt+oOBkD
2K/K68ZJsFRhLPLXZSSs13SuBGG/06wYM9+lsJ1W3s5EwN4Ux39lzOOAQFre1OgHIu589wKJmek5
PKcafShMaValVk/xlsWlN51oB/cQbW3cgVjIygeAt8JY6AOpS6RdLPKI2hgWfiNhpO7DDFrmcUri
S7tXBGyMOUKAgTvtVX98IRvH6XQMul7Q8poidu7OZuIxsD9+v4U+QKbflGSB+0S72Gak/hoef/po
ZH70M6APbgqGo2uBBfzT9KO+gdiXq02JOzfQVWZ/ZQZiJin1f9RMemCtsF5AO+XFO8HpxP+YPXZE
0LOp1gw5Tu8PPFxGFM2pmhJ1tvqiRowU/CbocXbcHnnpBBI3plibTpTDhqzuxRVq6T0y+MknkFQK
LPgnCmeyKon3+az+yQvqWt6VVY6Rd8wAumjEUjRbW8ayYTCTO3ZkP2MqTAcWckLwFkuAKYcT+HkF
IujDCXlGLTtlebCMVkFdmIssjWrGa0hA4aLzc2Z5z+GxLaYFre+8CgmdvJpWOA+Dh1GEf5CLSic2
zamKFsKI2e7taBHCUmVBliI7Aoi/x2zQh8SQkVRZCa/64oxywszMPMErKSUP0xNIyVYjn9n1aYc0
5fGt9JnwU/GHjfTgO3FtaxlKqi5SlSQwAERCdvki+NkfLbAJREFkVVX4q+C4c/hX8hQ93G5POSY3
k9nNCi2ZfZ7TAvhf2I2LYMmUsx+e+pm+d2ODNPdqL6YaOEGU1Fm++KtnwEsDkmX0jPHy3QkF4pyP
xNY9h8NqnmvIT0ytyLP0LT9zWnA+8HQkcxbQKmgN585rnAnHF0xxI5MembquhYERQlIunNf1WtsK
ydPLT6jBAH2j4mvOi7Hde0Bi5NSo/eMph6kDQtPxmOvQncUZv2g1loAOhi0NOuO042nIdXkyaBZD
fYQkGtJmlUs2mFYv1O5wXZ3Jb2KMMggapP5xteC80Hcv466sm9Pi45eC7xaat+5nbWsF3/Pug/49
9RIEKouYGzU+IC25WfMKVr7STFMOlSDIeohn771PYbQLqp6X0W+Su4MHRSpSRi/xclFSQbf1WFbn
1657f7fHEpFitAG6aEJhI5DdCIrLwHwVa8HkzT7Pf5qX5mG4KStrXbYOwr1wqUNB4PQ7n3T6cfHC
UeMeLoMIEvxpVsl3xLpziYXBeJos9wP4mU2MLFErL7xGNSmNLr0QpFASoK/XxCao4fD289o/guaw
Q4DxEO2k/cMl3PiQdWNpwUI2Kj8kJHFyr4yeWpWVjaLIgGvQKjiUFXhfpVHj/IV+j15M9+agi6e5
7l2/IcslCPVS5bc/VvujLb4p4QhYRbLML8KRsdw5GSiMjcRcfFtIA4G4SR4DSSPHgAQoC1/yt644
zaThmsOWGIZkCkVVeQFv1VxmP+k8JHTBTgBU8ifPBbzpcd3rnFPI22c7fHE4+8/e8R5Q46lZQ/eu
Gg4UQxjCTQ3GAw/G1NquESHqxNYMwyQFGBOM3qhupAnXMQhQqW14ujFS/y02fMAYuMppm/+MFNrU
OjiVg1mlEcSZexYtstvidGvk0vs6YVXlqS4jnthV+/CkdxaFIQWJXaPjPVOvcFhh5Q7squWB0vFr
EZztrIic9QYhhzEZtk2txC8GlKPMNHwczJx/mS16W1bfr8qZjNlZdvzSSu/rBb10AWH28VFQG2Oo
k558N3qYNHeNov160vZQ/sDHmmDX56Z39xVYDeAudrghSwtJQMpEQj2fNHCJ5qLu8/P0d2nrgFdb
MVoJqSDd8HeG0HAQ+iYYQsxTHLD6sR6BNQGw0adoPTYV5r+rBRbMxMadd7+ZyVyw+PfnbjgCqgtO
xsXDbQwJ9FEzlnKFN+Ub7/P3W2sfLySq8fNcDx7gGGmRWbP5Fvc1MXDJ6iHrWn2/NKcD+obhDLM3
VKbcyYBawmczc4wAR92zo3RiRfb4qbe4G8tZAWWaQ2XwU6cRKBIjFzCb6FmGhZW0mA/neNVwBqoI
mgw1eOp9OL3p1SAPn95NRxSGnwDkvhnAQ6aTCLgkMeF2gHSiF4AB2MFSkqxerCpxK2uA1KB4XC+n
HcWPvKweJbRuswsnBYJ1zOpEO6wmwBvopW3M6Ybg5zjm7sbxGMNJtjZfz8OGrrhCtzQc3Mhotu7g
JCH7S9M+MYZjhzalxY1QvTeJoLt2RM+iKJcDn5JPZT5ZOIlIWYPChrdQjltMQNT5xinyLO9MmibG
/0/k82o5lwJIeZ7L4mw/om/l/nX/g4Dd/Zr3WXeDcKcddjQ62NC9hC9gRewuAAuJ8oF1RyP9vikt
NmT1gk1pintHXvYw8T1xkE7Du4bm3dTqY593Hi1jcJLa8bWvyjil7gadylqNP/I2JhMR5zTQ9o9x
xYXRA3/30CzSjv/8+OTIy/X6DW3uS97m9psWfzKDgi/ZGU9t6FyWb2zUHJ6IK/yREkfWYNuTdtJM
HC3abgiE+30Ip+XP2PD4aKf5Ov3rwLB23vvhOW43QQVFV9clCCosP+4hgSJZh7EnBpdFYmIeVleH
girSaEeVqQKoSG/7jU+12EqqNipALuslG72aRWaq3KWRsxN/ygpRvOjaWg8ArE+SfcMSIcvSI9DK
UF92OnSMPIFwYbBYhsFnLkxBdVpq8k6T8fXXR7YEgmgeJVBYI9ahoeydMj7UqgnzZx64a9AbgSRO
l2Y2DcANdfzHIO+pBjA1aThiA/Pankfrcz97HbOz54fEqksmJMS6PpP+n9+7ijD5JMPUO4tvAKbB
shN/ioglWdQc4YwENE7WKG/OxDBmqX/yflbnHyOyVVjoYircVG6Abz/Q5m/75d7AnjMLiwhBO78x
qJifgIolNih+/DNM/YEEd1t1/8q9QnoloeRUYXjtPmsFDhWl1JDSOuhG3HkU2SGxhM0w8twLZuOd
N3mUccg1oxPy+T3eFaKyijt4au1YMMwv6Q65DeweAYIAWLSc7/5IUHeWLDwYYmVlqWyGoARwEasB
4GBtSFecx5LS6A9fY2uKneAZAgM5CDi91mcqTgMH7xSG4x9kzAnvTMRHbKZb4stoRKpSvg16V4ek
teQrwJEiK1BSddw4TSn+twA9zrM58d2SkGI5zgVdNsy0ICVEl6QBYesqkVZ/tqvCMG8xuB3P9nfB
x0PwMBPQBMzf86Jcq2o8ett77xA+LSmIsoxu1QGxRWsgdSSOWtxkdnvod1f5yn8XKA7oF+pTowTq
zfcG7CEnZzL/OMkylCwsxbaggf8gSEHJHH6waWkQbtK3kCLVycKs4WlTkqWVvLQERe9XcXvZap3l
YMILYFQZyQ3lulYeCEW1ChYVvAwN1du/Z/dCkCmwGTJTxbkbduzKVnbLdoY9hKoeFoeX4Ntu390E
iPOqzM+QW132lYprytZrYsKNpTSWVQTA8CUHqYrtQVn/zDAQ8FudzXxsleMRtzC06ThgMGsqsVY5
mAVSlDHF63eMfAit72G4kjxnYLzcRRvxJhsOgE1Xh0xA5hT6pvb5bGq0/IVMZKQvN7y9hVaxezxq
VnK3RwaZk0qQbIMCEQQza1EAtAHRut9FQUInwj/linN98JwtQGGRk4HIwY8O6rfEXaMMTPoeDE2g
WSQyYuDmjHtsWyLwGwGsKFJZ/Ix19pQ9O0+OYcPOjMAOvgUL8fXuP2VYb9Zc5nIYz9OVf2I1BiwR
CHmfN8I0Nb+1f/b4YPypOmvP0ikA9HHEYSPTwE0MWw9kGfy7t0gKDHU9s2nDrMEZ4/9q2OQKhq9c
n8arKEuwKgxTBUp4FiD7DaJolobhP5ZxQOUDNkZHvFFKKzQrlXCCG928Tx5nuZ8gBCV8eoUWX8rr
GsgwtMzITC39HT1CgE+aZ8WP1MEAB4iGfichoT9ziCz8ZFP8+x9Mf52/M9Y5Nnbw/u5qoWZy7Qry
juSATXrXLbhFF8LIrOi+Hyo5Yrt2BqcFNu1ZtCRrGMcy+9ISH2bVldfCUsnumKgfahILRR7VsrqW
QU/1AaPA4XaZuKA35apwnJQe9co3QoLvywljXgrrvG8lyAbIA3vxO7B50SN72mIZTjON4/1QjBqd
MGk0tCDGON7/n2+uedLHQVQHVR2GyFe8nSqRTWlxPslU1raYtomYWslHrSVNcHE2XipJIvW/LZxf
EmJvwTwqCE+ekMQYbqi0nsM0F++juWqFTmJiaSBL5e3MTWrkhdKNL1cRSBES6oRg6JYG0SMdlrBu
BebAp2brj/Vltl3lZLHIQf83xM2S8RtKtlWrkF7XYoLtI86/Q22Odzyn7pHNjet6LlVqr0Tp30Qq
nOBr0UwYInya5jU7IOlkaWHSQ5cXVFtT3Zzy1nmR/UY2jHn06+z7rN9go2HftRu1vcSdEQ0n+0tD
8YXnwnTwbf9tglnx9jndF+cfAqbMcYp2zp3JVIpzoc4w7qOMMpDgYjh2+UA1iSj9dIzXZRHst81g
2sJ7QuUhKZqiWCXEr54XqUbi/LMa1ow8faos0Et+/tERFtPpraD/JnwY51cJGzmem/GAf8hm9MwP
96ZRLFapRrXnXA3bS7GiYPuBx3c5ble4Uk/LP2KFfrhMUAGQgYQ3VdUyLxoBIjFQdSfxOVpJWEhR
8vCAhYgmSUSRBaV1XwaLSSGxLj5FzzYw2nFMwsnAS4Lb7XVnCPgWWWxc/ef6WBtkACrogjeoyGIb
mbV2LEzFqaRK1Nd1x1HhSqVV6lRMEXNQi8pN/SD6nRAbu8+1y89vNg6Rd0emyw/iVn47inRiFpr0
08gAAvfMxdGoHX1mKnFo9vJdxNkzfthdOBnjNnA2fy5s6MaplBPbn6DrorxdJclgELdeB73JTLaU
AlZfaG2uNHbJaE4G0xh0W9TnkcM9nSg8vF4eocpmcmGayDKEIAb8cSiUUFk6Q0ITf/cbEml2JFxT
ZGjliW5BrCrOHv038QcuJljlmuqYqd0ubdEvxAKtwmCYaHf58wT3FHd0BtCbk7DtCH4x0U4mkKts
bmDK6r5waA8YLp7Bezwi0QCGyoJAV2duN7fLKitQC8Lha0R8QyjNwEGf4Ic7EaCLmInTXoEZPWf/
NgtqiaqfIaltiqOU8kYkgSNJcEE/PmMJU0HbwSc21uygMCz//rIiprRlFsp+uG8dvz0khuU1mKjj
5ktbMboHihuNsIbsreQqcNjMxe6PIgjp3H3bibl80Mlg1TOiy9k2QeRoQiwVwo5Y+SRlAUn4XR3N
3LGpbHWha4aBhrmpmAlClKpMtf2fxkqToiDONuV/brwoMSLh/bXpL9yN6CAWGLleZc4CdohskPax
FkIXov+t28IbsISZulWUSoAMBYtxAkRXvnEqFzGbgmTWccOGJEp11ZCdXalXbpnjhpdSEBp0QJwq
INDccrVCVDYpIi+bJIrB1tLgMrB4zAIc5C6f2F9xXglMVfn0+Yh5u4tfrk0CgOdkp1Sp4H9omz44
eero9HS3cmhRKHO3j+XUxGhhyIMl/gNrSWAyCxc7c4sel1yzlbO5KSwQrPhEWiSYDv73kDjLHZ15
iqLdLqRkjtN5y5VcXvI2Bb8lERPbAizUpg0KlAYyql+mEqQBqpqSyLI3K+PeIVlt3JM3+sfbAL8/
EQ8bsm+D7ZnjMCglNo/Ib3nF2kHknmF0NVUTS9ZsMPBIafj1xSbIXZCz8quZBNDp1yo8aXM5m8vX
AKVquNoTSVUTg+fx+MSCPuNUCpI9PfszAjgy3nfOerTn7eywdb7V6Ns/ZixXgmV9IcFADAQK3fgV
tItMfXnEGG8dvBK4VO9wmc9FlefM3SzNRUPFxpq41ndmC20cNXjx/Fld13Sqwcq2ABD8RQ1mogkb
K2hfIvKUvaNEdJqBicF070biid4qvoD8Tu5kSlAm0rQPfuVaCA700cIrcFmb+ttGnsh2g+hqb+R0
5JFnn7u0aKCUJy247OATqduea8gErKgSYasFLZbUAYXzXXpHP7tna31L9hM2zIdZCVjslk2ecpB5
Vq2GNX9nv3ifIynXO94iOFpI+0CscHKW5zIwzKt+9RLtyDqxYJoDDjzsWaJOGJfwWKoVOwr/Z7LC
z10ERoppH5yQI0ABDmbv+Q1T7TEB01lJHETxpKbriBg/aH3axn3UlhQB8NbeI9TC8xTAfH2r1o3M
Fh0B09WrgmBd4lKOzUcqoHZDYiOqNnlOELhnfYt6qdaEo7MpC39BWev51dWdMFGuq2j5wXSy0fiM
wMZpXRCStXSt1lqwrrPm6fgIzpUFvUb9Pg8xZEnceUH8tRZdsdDHKkrU4nMOwCYZcVviKKZ6uABa
9s5nHRJ0lfC3qndhXKvzDGw9nvNUvJSfYlRVM61ntJfyPahtnM7Q32vfLbSOVdT7l4JLHHpj8ujH
8HEijKxuOO6SsuFA79SWsqhE0F5ROuRle9Rh2Vl96UYuYQH2OSnq0xY72PP9661qFmZ4SSptsvr+
dvlhM2MLcEYo9WHOQBkj0l7FqXZCFtMA3SqqQ/2i4wBLnoQxhkot8npI1zUiwnMf5oNf0VisxyBU
kiMdRBz0KjbknoZQZ/8DlDwDR0+QD8WFQIo2zDosksnZgJqYDWHN+e+AN/JEVZbHmi8iiMrnfJ8s
VxLTTHfr2Zkw90F9h350Egf8Pw5GtrKhUHYn9x8eJL+NllNXXlsmxjpF3bPinMTIYtj3AH9ar0Zz
eZdPFhGUzfL7Srt9CcQPeu/gNQng+ZewFHUOzcumUuokwZYZNHI4WJCszKRDvF6ZTqJD2FESSlks
R/LYhh7YIS+LFtJ0CQnC00mIWbL1vMPQijjF80S0//FGn/oREkVA0bsgX3tM5CB/cI+foZ+oK4r3
o2HZ/tl1Z6PVdNQkPjIaW2f7pNrCx3dywvPX2cw3kSIkIAHmGEn/92J5Y258RGf14etup7eowasW
VfKbB0iMl/PO9D1wYq364v9Wt/JfC2b3k1e88qNCuAJD0zUheWWz70YwFlEL3hLytFqL8sZ3N4ww
ZLB/agg8NkIziiYPvnWpZLhMf+gDZytq0zGCImWCimaxihowpAywOfGfGq23gAWoJafwPDqWJ06m
C6/AKnFCZ9/1DfHEX3Cbw9BhR/G3zakT+ZNoOlmTiNBrksqHiTEFStqE2cIe/siTaTXc8VArfT0U
gcfBBv5DFHa5Eni0zrDoFP9wwXSDTOTBrFSIBq9aMz/YKiWqXQog+Npw/LtZ2ZnVIrpZ1IHnZ/cZ
LFl8ATm5ZjQ0oGQpTCDQo1wRnhXwTplmZFh7JpQ4fJ4K+1WJxLASyILNyoksyyj6X3Ma5sauBA0e
X2srYLd16OvdRj2EKd9svv84VIDB08Ypq0paUEqHtdBF2F8QXXv8+N8tr/2SUjr6c3HAgmwkutFz
4U4qcP8/WqSQiplnWd/vkHJb05d90MuQQoHe9e/HRoBoaJClMaVNCiW/NgnqKBnImufkzKcuzZsN
TOr83yxNMzh6j/P9vVTrZ771Y1Vjn3+2n0cFvXrNnPerW9/7dFENQAcMwsUftGIY5ADJNFJ4XWDQ
cHaeO43p4+knzcXamb0k2GTo2SJnKWoTl/8+wR8AqZbEG+PPC27C+fyYcd6irpllpmWyMekbLhES
gkbB75oyuylgHl3LF+0pX7pAVx108MN3FMZfgYCve0czg5TXVxyZwXbuxME2Oz1nNn8gnt0HZpoU
/uqi4oOIB30/6THT4LspJVkcAlVydEqsW1pLjteVOMGYJMnJubMQJmbMeF3ljQMCc6RzDqFBL79z
mqYPOiblHzLjUu93NWdtUrN0x/zUTeNUFiEkNOu5qtC0uXLIAxACBODk8rK+QtEy3OQpyKUng4je
rH4a7WaozWkv7Gk0UCJp6oFjDPBNTiNdqA2RMtdiwhUbz9wToxDVhk8SumnBc9Nb+RP4TvzEtQ7k
fVE7n9B89y8mmOvBsqGaxOzS+//ly9Ji6VsoNeLjtRd3uSlTeNQeueW8EbC3EAClNCXCEX9eb0ic
M79kE2fwAjKLuxagb/c2Wf2RVMQMLpLFqbvhr/EJ2xEwl8G4/Jz4//VUiXjAogIPQQGpOH1xdqwc
8sRjd1UxAQWkgTbY/6ZRnzdBf8hpr8ex6ViyaHa05HGxTcI437Y3YDdW1hUzU13hsRfFF1uiBAh9
UenfNRmXxxXQrApwr/kI7opDNxhoBs63TrlxB6cfy99d4e0su5CkIBPf9hq1Im3f9aKDSBba5elu
c1cW6quZX9vEiDAOro/0yK7bMRM2bq8rVqOPxLFm4TuEbu63p4H4k0uZmEvIvCGlVJb5sQkKR3Xx
4SOfDzPaACHa7xGW3bNbXZn0bjanqLGVqJh88dClDlPuTy/38axPRr2D8sVE1+eA38ewgX/RPPJy
CGldnrEgBq9/sfHwqauy+0ObSAZeGLbTkUgUgj0SSgN12S6wnXN+9oipKsdbatz2KvEhbjUwHlIT
CKG6HA+rmKcRRoYckwpf5iKO69EPZfOJp2GLP5+EE644tkKaviAUilsZk9tj2k6GHTKb3a3HDpyh
CFekB0a7KgFzVgyukglZfYq+evYtCQfW/F02tyof1SYwPGVDQjg1MiQQkpccEknz/ArH+7yLtLKw
AxqrQmNGJHPlULZLtGYa0BHfD17rnMabNPpmpRzPmP0AQoOzpnLO1ZZ72bgVLWUkucis/NFF1j0L
2FMjS44DkrO+5Y+YpxxVg5ImZHnHQ1JH3gvhiN6lPYptXDPEHpqxsVbQXNOQT5RfFbst7q7IL4YA
jRlqWG2PF4qT60l5vmVCqm04Q0FiTHjbxLS26v1PvpdaV02Hc8M9wWWw3HZKQv/Sf6Uf9WjGKuc/
nt49PfTO/723gpuZPzTLQNwNC1FNZd+k1c+CyevCwQi513yz/hWG5LiBl5Sj6wAPktoe9O5sS05K
DB3R88khGBIBsf4EUox95BakGN/DfU6ohAA8C9HidEqDpODMCvyu+788grylaezrvgvEw36H2Wk+
2Q12lcDM8R1UuC90lYWrAlGrLNbzJZACAVllPWyzy+uYv2ZrcLY6uch1zQ5NO4HNVeTCO48/k3RN
1uuYVcxGfv7fSPr1wrRAws8nnqTvv63Ln0jev9vQPDuhrQVeRjhKXeAVwNiiiO31bgvqAKfGiWJr
bipQgaO5QiFJHi+nwiURo4oGki9ssSy92PAVU7xga1Td7HF04S24eJj+yuTIv8XQM+PmogBwvHxw
Cz4MC0CiO7UL0LqSRCheb7D9iw9Pb27o+NPqU9vJfVen2zdyNBweBwiJx5k26jt5zhe3K45VfNdF
D19zTyVo5UTd3NlAENci42I00gKl+p/y9ekviMLYZpWZuBi66t2SB03q2LXm6nUoAOSMCv8385Ui
eX3KnJrs1kh/ZTzX/uXDgTv/5wxZCkqJxNWELCFC5t0+8P1WbEgJ0U+X4qjpse5Uj/l+siPeL+6A
HJuEW3t6i5HFkEysT1HrKaPUVfR80hcFbYvEj/glUUpGdkDesrg+JQfmkgxlh5YXAP1eFt71y8cB
zB1EsLaoDuAdXRQx8B1AHiBbFpEq82iqr/D3RaiAk05FnGK+KhDga4rq7r1tExAg7JDTQZjGEevg
Rrl2C7dEEFyTteiB08NTEf7Otj072EI46C0MHeSJu3kd5H+FME47cpuSJrOHVqnwjFFhA7L8gM9k
8rWjto9Qk4mPzhowwXgdG27N1mLZTysoC1SshFXFYyn9DUPKJzkrVytGNItss48mQWtTa3v6st0s
/w8vdS1hsYHD4Xjb0XI4jxAxY/jo9iXhrxzJcTOt4u3ezCaL0XlckaHTSqzmf4RMh5fsr2vuAxZI
W71NuxRvi1cMGVQnoOFWSGtGEdabiHRV11NF+fQDTI1/RxAx2P/LQ3n5Cwm1ndKMRERk+9fij8SU
IHQolTDfwr3u95zucPXLeTGp1GOgy35WSkT7YdbOKsTWGIVZSG9QkUH00+/PRGKv4fRCx1YJLOu6
8HKNGT8UDQs3Jv+5EH/byEhqWMsC0UM6gTssc/VMv8sbCSnlYybEFUHOFyahAf59EQcrRpO4AjfA
LP0v7LIa/M4x7cwb9enENRI1OiiLT831DWoA93DSdcihzi5RfxqH4DtBxD9n/iS0ii6VxE2K7RD2
uIUPYhAweDm9XwIgjv4eQ+KAArse0LgXHfTtz6zk0k29RyiPXNujThBNsiRhQMSGEQfieLw3pGSr
+fYUjhKEe8h3GxxUdKvNL5HaAKr1LodKwUPQgeI2T4A2CgQVeSytx7CioKUUREtPtke0KL4mmD0i
DSp+VWV1qMky985ujqqLheRNIElV2eMJeJwWu65Edynu3gUdztDeP5Wzb6OiSuNQy9/lhbqtJ294
SW6LT64e7S7LOLSy/PhO2WFhoGy0h49uR8iH72GCwbsKNsLcxhyHlu26pvjLsfuPuorA0i+Fd7Cl
x93zjGzSr752gblu/oGWuboHaG7EsGQbwVKy7ne63LoOrFjG15IfYh8qAOANN67/jf7DygiungrX
PqhrJl/rZVax9/MB0mRR1HEFfsqYUGaqIWCiJ2VjqsDujAcF4zxsoHh4CUG+UNR52QgukYjoFiVq
sk2/Sz1nRi822Bpt5w3stiDbnBRaaZjGsF59c/OhAB9w8ScCtvS7BBcbmvTEGiNma7ciNEdTjGYU
3q5UOjoZfS37YXFfCJWqGBk19RTlHGVYezUUh+7RvPg3mKDmlrd6CG4p/Njr/0RxhiZFJs72gDJu
iPv6IIURBHGjIMtlBjmir5zVl90dND23Ge2jlIxcNV04WxfQPjHzcnbsquaQ35twu09Y9mtecggk
6UxytrQsXzYYNz1K0W1rcoPlqtVSIENpK0pCsezN2L+PR1x6Et59Y7tbhEt7oGGn6TTyB5EeNtxw
yEWnCd+egIy8yHcPJZaSHgl8Obe3iCB8ta5RTHLXRuCfbZaI/nJBoujQg2XsON3Vt3HbRyl6ylvB
be3EGL5m2F6qNpE9sfR+xoNcrL1B3kbOTNFWh+ftEBdExFxN4Nja6GAJDqJc8JxkeQ594ZEgm9J6
MscvC0Z5ChUFtyvpv2FUTwRGo2JcJjW45mPTA2IaFdwko1E4kc0dwTuXOmN373s6UU8Mc8dPocg2
vMcnO+fKVcSa2VJ7zcwvPthhLn0m91mnZP67jz8X+n0j3KhHLDTnEhKSpYgwW6OCfXgb0WB7LFP4
qEHZ3co4oa1THUcPkbTQAI01nTlzROsQZhB01iaf1HKiFHRD+p+An4gK/FR4h7iu4dg8jMOmxp/3
K/90v9NcwwyvGeWlsRf06CLh/3AEi4poqL5gHvVgk4S1C57wmf/asfyom20o51tl2bCSceGON8Il
orRXaoKY78/2JPkYNH7W1fxpJDVK1cF0yU7liYBqtH5bXiHgW/+x9Z795F22Wirl65GeOlQOTo7i
Lh8LQEGKlzEdKbwJrK5VGmQoCQg5EUWxxD8L6T/JQN7zq+JrwRwSNgW5ASdAP5BVgUyJZBAtoy2K
JP0AtxpWjstJcFdwU4g5u09JCpOVR7goYnei6vXDNK8TEq70UKNvfUZ8l4+uSlwI36hQ1yYQqOxz
wLvBl9lPc4QOu2UOizOlQbNAxhRsZLMxm1K4o68a04fZf/6yLven7U+aUejryMBE3JV6tfkIpFme
4+MtnEhueY0wV8hk5fw1wQcaE2ac0BG+a4khBLC/NMwOYxOROgyt/UwWTyKuKSMDVBUEuuln17Vi
+KY8BjpSlMWeo8NIQHDTzKUb/uHnLXmKOKqRjnjwmYzQpTbvubci7Axrt29XE9VqaO/hI7WJho/R
Po8pbtkwVOBCWyJYfGkz9Z3cEqSHt4IELJh0BETAEN+8X+/hPvLJxc5QY0jJBl2aAWMXmvVk4nvB
TYbe8YHsG/42bcqZAIv+qLWOlOujnStvOs8eLTKp3DW2FpkxiqpZUj9TKOspdCW90rlkkLuVdP3F
+gfm8RX//WhLNGid91JppIEDcdzWaCEB4HmhbRfADL0c/0pSKq5/3W/AWxHzTQhc5u5jhY99ixXr
v/yeFqtfx741OTy9+ihzIu6Yc/iFLVYeF2AaKKzCZoYCxpI3/8yeIKCX6WyWTtyrPCYm9ttspfG+
w8sjMGINvI18awAyOqldGvTsrQUpD4t0sQFTu9F1MqX4mI4+lESTQ5NBUZfV2MJrF2Z3Pt65KiK0
D+oYdCEhxn5GP+6VO25JkgFqM2J9sFbN9Nw998gqSobb2aZer5imJ1MJEPPneJR8DA3Xo0FdLvZo
xmPdUCP56cr8Ue5/j7UbSBkfkb+kd/ttBunc1JrR6Cg4+D9hZIKt5fEIiATcnE7YRKkkdAZQvtdV
lAlydiAGRyUrBXEgSdea3cCjZkCVCtXe343Kmbv4VIsiZClIZO2iMoZyRigqy+ayoLUHy9MwdftH
uQQEAzrQN+Q7xsgtAJE+8hLgwxU3P8p3AaOK6w3n2oF/iFuMlAXfRWTJ9eVETe+B9ISd/Df0wJBI
YzJLgxsbCiX+gDlDRwWDkTK0cgHrVhIl49zp3TdW9aSuUJbrTTY2Bxv0pdG2aOwqRfX6xbHm41+W
UgACUv9rZzDwATbIoqaV4VSidstdg42tsVt74SG87E0VdQzOUNXqZuuUm/J86WZ7hTTBU/u+xnA7
hLPbSAWYtPzx3q72ESL0AQYD4L07YXErvRVXJ8vob7nOfK56LGqI9ibFiS4vDWWuJw2TRZl0QUnr
vyeFdZ+I8SnWYS/R5vYCUuQ5VMkqZbebdPvjFixeCJcFS77/GiNlgZFQEww6LvweXX3EnqxffYJn
iKRX1kWJKapjmaWYNumbzDDPA9ls0GnwbhufHvRY38a3U1+qlOee5Qmp6eAr4LlwtL5MRsEWd9GH
E8PJhYuAX+o53Av9Q3mkuTETaV2xFfrt3sg9+kbcJ7aZW0T2M/GpBovWI5ybF2K1rnwIS/l/Vj3N
5yRL2HzLrhzj+nCwMSIfHbVbRuN9udhmT+Y0s8D72L6FwTLxDkqcQ5G6O6FYN45KrwqTh7Rp7N8j
va6TqZ3SJzQqYfOjYDeR9QOhtri8ndrCwU+sLgcdocCingzQo5T9OkNjOT1JtIhxLsdNAd7r1loD
kxOsxbHMsFUI/O8FikXT92EKGlozEA92mee5QnBW8ogKhbT1eEHLDsUUZ7M+e5sPHpkrZg5mm2yT
AWpgW/2RWv5Q+4POdRw/WgRtPpfLp8HFR2hMgVei/ZS7iPbsxaLJRv5ExCeZdr/rvzD5jcKn74nO
72LsRTQ3EunJKhYX4xZC61wqOEW6TwkSb1yAb+ZOvPrncPJ3bZT9bnWoBcTLpy86I3tVcbwMeuVv
1gwt2iF8pcK7NZr6ZmWW9QL22MVhZprTznxuRB/X4c/aELzVoAhYA8RXwG+1YGcOmH+5kczR6cy/
HQxfdctw7lzHK74vDY/9PV9EqTq6JV0G0TLvqYB+GBOhiTOOPRiVZvndP/rRFTbS4Xec1yQXuF5i
LWpkQ96qiskw/9LmNrYEmx/bgsbjNw63RVSe4beBz8WmfmeBUOTBpAGiQmo7Ziiq3qr3bcG3LE4E
F9iOvsk1cQeEiWYDi/8k3+GCO4x/XgC9Qur8xa/N77+ecnh1jL13cv9jRtTIN3TDdVNAn2CEPB3Y
SZOKjiy45Lszi5ZwWEbcyH7qIF5ppCwC7xxDTPG5/TGaJ7wdVbnhzF4c1Al65/Kc7V2KZ7lCiHAq
TyHGYcTwlkEwZNJGtiY1I96RvLRR6OlYEkJF9I6IXaBSZYZFT3d4K867k9mU846u3ZGo4E1eWXz7
Hdfp8t8wp5UKyyJcuzHsjLaWwHCZZP11+a59Z61NdLOH3Nm7+myprhlsEaZvSmJVFpZRF5GpAUXx
L1hMM5U06vSX+pU+OF/tO78c970Sb+nWqy1Q7vAYIgRv2V1nuBEX900R/fK6dMG7xMUp9sd3yyWZ
U0ftlethFwXYd6tB6p566/QfgzHFR7V97F0NOdqkTZF2MPDxCWWGRuxnRp4QCmXmc5QNUDlNYqCt
8vzrWqFkDj0GzrvjJJ7q3aRAMGxY/jNB5LUpKAQjpA3nE1TSOnDlL5zryUPRUITPVOGZE8nlmXcp
4WdhfVBVslucTFs3KaSyAglPTlEsojHf5k+lYvp/5zUY4V74sdBVtcZAB4Ex4/7Dqk7v/OkGkisZ
IHx9j2EErGOqaIAUDmRE/16nNdfUx/8QBOKUC8Gbll67ZvXYgLKnAZyz5L8gKbnsjtPXqEIXXB36
6xOBRaVbsgnVqKB7H7GUm9XySCx+WzWD4+vFuMMMeK9z+3Js92nStZyHeSVPRVF7BjpIWtD+VYF3
ELvIM/XYJFZc0oPhVeBLWS97EWU5lwoX++dSSG9tL3YVOWWKocuz5LuL7g9GaX2cMVbGmk/CEDQD
XW1ZoKm+wNM3K17Iy2To82DTPXwOIqJcbTHa4mea8Br2DPuO/mmrDn+q6dzmO8m5k6PaC4XvRvMo
vHZvxp3g5OtK5HRMHMVhx7Y8NQGnysULcjFL7JMwM3hy1s14Tiy+GNFOPtxSJPsOT4koYRyA4/wg
lHcF183Sic2SRyQ8mVTKM7KSyvSI0vJtg9KovPsf2VEk9yBOji7o4N8c9qm5XOfUMxCltUtvKuM6
NvsJ1n2WbLCak20lR9pJWK78z79CtP9k4mgdpYfXWVg3S46laeOC+QzD+aV8CmmkITWbsBLEIOdt
zqAIUBXZ/hF0orhphZEu4XyORSfhwQw/3iFKZLVCqDTLXafniPD3PqHKcDKaMPjgtA475RFZrzjm
EqMh+ce7BQSyUDM0rQA/6ByEnXaYJnpk3yuzHF6UAB/Nu8F9NCEbdSUYkeZyWa/qSMuS9d5rTN8A
6aBHeA0PcJrr1YcVMj7eobM9vy2A/0rCxU9/E5pO5wCjERlwr0offQi62eoPl0T/5f1WL1p8J2IN
gEnwzM+W3WIJ+y/QbiN/j8DKCOkGOyFIVDxBlN1569ndfKH2YqWyXfs6BXE66sbx7vWL6JRyYASc
L3g/xOY31blD3/9xseRt7EN39f7Muo8CcxkT7EPe5GbsE3hxTh+bXQ9MSsxdhAV4znx8FEojO83Y
2lAyWtbWYhXYNx9p9Zl/224kJvp5HDmfVVCTK2qLa+3h1PTkm8YRwKggdreWPVoDNKi4SuLwav9n
3bBUxFtlDHJxrq/Pc9vnDbR8HRJ96VfxhBljDI7VBnyfhBAqfwmZbr4SHwEaebavbIGFNKJ/qPvD
RatnJLTkUqIqDOH5Qh5rTi1ZmJU1oE6PxRgZYYoi52B01U4hOTXChSxTzgxBGfoETObuu5VhpBPm
IU49tJsK8aekccCt9iuTsHcApi42HLV3LpACnzIvEZT5o1VJesgd2IQntvSTbOhZG2liwwZnsAhP
bx+tnE2+9KM0N3CZKIEJi72p8oEbu4a89ig3TSBZBAtVksq7O7Ot+Drthaf8gYabitcW71NwXy5F
pcoLoH0BBJ/m2rDwYhH4rlTyAHt9bpwp6LBCytD4xmmAtskeCiYjVnanSLacrLpeXTk3VD+hZJYE
aCwug9XcWVFZsqFNaB6V9wqVcnxScbiFx+0qX6JvTn33aLwjBzMWzve1MVA+QJMnMWHPk2hthjlr
ru/TYi1fLxuESlmZ1bdd4oKKQWbqcjOdVpndeoIf8l77fiFGqZuyihLCxsFgImYTTRmYR3Og0gE9
3OVZNQf2BDpz4j17+uCcZxdsCkldrmSNsDnwRe+j2i6mbjQEH/PmlfD4tFmoHqnw2vMO/irq8/k5
3l9M27aODz5o9/ebaVOjWJ6tV8qbP9oFD1gIPytpMEVBYBiHMQEVr8KqVq+SUa9zflbzcTW4n4Qz
p6PEdS8QKrIsPlu555MgDkV6Cu8q9E/6R7H3BoOLkm32eup72LzRlU9nc4Lgw7FoF3hlXSHm+2nY
lfy62d7y7mkg7Gy9jHf3durMuHnL3nLEd/ymKd9Gf4FFdOZo+dBrRqD7cDS52YyjwAXbMSW1cDM1
uG6MHvheKcKB7e/w8dXpE4LIsvscDMK1zgD8FAyDbm+XCxlofR/Wm7OwURYkxIGgtBAvq7EndwNM
ZD5b7DJagm8h+SQGTjJoVnU3LhdA+6Au8oDDJRG2rz8LcFC8rJg1KlVNonVdgRMdrx0n9YhizgJD
fHcqDfOTkrCxldj10zz7jxeuYiJpo6YhkFJLqYegVC6mSSNZN+82vXInDiGcTXgZmIzPJc8tr3AX
FwqKwUlX0n+uN6GuIAuFpRBFGFZ/uyame4f7bMEMOnL7uk7H0+eEN155td6BmaMH6f9T/Sxy6BuI
f2lk+JvM+LsdqaVMB1T+g2hbm96AOL99JGwb4ON3NR90blGTrVFkkRlpjuLaCydw5sl/Kbt15I76
cG/f7ooaTIfVYHvg6UEt7qUDck5zbHDB4d1sxIS6cGEstaAKCt7Jy5JWH2XaVFl96om+2Znn7yHD
RHpMrjK4NfmCafSw4SP8iigWSHZ5118+u4RkbB2VG9vmgF/T218cFD6e0mgy7JhImRKsDqJesZ7+
17b0jIzhORRABK3jRRG2uP9As7jPDqhedfGGtPSmH4hbfehzZJ/ySkkUUNRBWxes8EmgAqKHSfc/
jqGQlZ9TM35gsL6vxhPpg72pUdNNajqJ6c0XsoGqNxWBzZWSwlBz5sX3F2LhFYw0PW+eRZfGiHdQ
vytaGkBodyeRTDUgIkvwBu0xR3eJxj0MG5WMtomg4U7PajZ93neBWVkZh9TzDG240FebccewmqwO
5MrpyQqLCAY5iZ6b+WAL9xnTkM2FJZT8ppYHC0ByTQv0Hs5Fu+rYT+Vg2ZTgZR1mcdf6Re63sgRV
6uKopYqFThmUulWcqBFjvXqtm+UOCwZXM/SK921UwJgcAZDHnew4bE2Hxu6GNuozmqM1cdifLe9S
12jjx/69eTUU3ntqDsDRfGESpl9YqOIv929A9tq8t6ulCw+f4S+GIK5n8eaPG5t4U6kNnmp7r5Hw
hsw0PYLGCC+7ZZ1GSwsMaoiZDYKRc++4IMkstJlpodXseOVcGnKg9BYSsY8uilNWFcxEvfKoEoUN
s6jPxNpXQcofOV6Lz9B6+h2JsX1Q1aga4I4trZX/XXGdsPXZQLnH7uorKLJWDW6FjCF/7DUrSk8h
/4RbVfLYUAY787EqH5Enbke0o6s7dX3JTzsH5RmezJggVVqKqyKFR+AqamVW/vT8idg02kNOFxTv
6DdSx/v4e9zvDXb2ivSC96ZdZkL7/sW2s+G4d5syhoF5Sm3a6ahJPyUPSel9iSCEPs16gj2kCfQr
pfX+DYbAynccaYFZ6BO6yPxtyXl4V/zutdrGcSXM3x0jRVZqpA1S6Nl4T2jRNaetFeloSYT1ewb4
eVcYEo8rBb3FERKf/1CSTECxl5+5HynKIOJlt37yamyt21ndeyGdnyOJMeImQ30dubhJXGcC05UB
H94SAYOWdUi1dQJK8WAnHGXR/ij0n6uZwjsH+9FatgDDhRQLclSFVLyoOjdkozL8At6e+EP4rUnZ
1Wd2hvpRXmVriTJuArX1/edkSE/CF5N1dsnS7uDSjQoBkul2mYcS2QLcXKNE0vAfC7eJH6WG0Bqm
dVUpH6Hjuov9Fo1rqQnkIc8hSO1h23iORaEtJJKjiJwJ1TuEB4oiloGj5pr00eN1IqOolKCfzGGe
j0gOxezBGC7ZEbObGmr5xMNmWRHJnbnsYyh2i5Gx0fABTHxtmC9W9OSYnt24eOcxVQqGqaPQtHXg
tjS+x9dUa83Q8TEQGu8qsBQzgRoaDL55gO8O5Uua01UFa8QvOmnkDRAQI2EgrWkhWDsGPGLM0DLM
YfFzFp/CMxN+wYxYkJcG8ijPZYJLZwhzzdOfWpWcaXIaNr4reT0TqoOBaej/lYNI+jTndiifru7S
YB1W/17zH0yRKMzGNNfCS3fSUnX1Mpv7Uk5ddBKqgiso6zchRUbUvQNAiJekaFw/z6kHAMfcQNQq
JYL7Ok+qwGrpvuJyfnbYJdtF6zdSTWPg1l3QDeak5N4zwSG0/uVQQTGQNjCGzaCND9RNVcKqLlWy
hoPWNswcY7IG9x+06lk/j4DHtVSvlfz/Q+1ilsagYwDsK+sEu4EwlIUGPwL02BRgxwbIZk8w6FD2
aNniv/5YACbc7i2QV+fceRnzZy/bqB+1+m3gGkWCUV6BtEf8ZJFLaUyOd+hTGYPJThylhf6SZErc
PsDbaNkoyhgAak/xNXkcyfu1I7r64cHxj7TE65aHW+0Clu1pU1UxHubV238G9niJOJEdEi9blw94
iuLWyE9L0DhPtFOwZ/NUr6oq+/tbA3VwHTPJVoGH1IsRgxBiTrqLr9GHFwXL3bWuJvXaxLA/dZxo
ZRs2wKmDbSBzskhnqGg8pZXV9LrCVK2YSDclJhVNNX9Ep/o7McIklYkyd9Axe4jsG35i1zR2B/fQ
ldPry4BzcmahrxHzVapJxSe6N4z+ZEqXf7x7Qdu9DBbD+rm06jDAAeoA9v68A1xtHP30mt0xFlq3
1BlxeG92xcoFIjcaUNQijEL4rcU6x2Oz1U1FPum81JxPGy6FsqceHAgGQDkMQRXlqoFuXlk6CEc9
stz86V3C8q62BkyOwfVkrjHrDMBvIZdts8Mpb9gD6v0Ijp94gmlKN/khf1K9+fr7TzCk3foZH4Sc
MBrom1aDJs8BKS1tZQT7Ky5sEl1T5Eqj/puEbD7ErJVbPSXvu8QenoO6nBcur2o8uFmbHRwii64s
f2qjHAjCVHp/zf0arTDroaN/NaVDca/xjCsqlpozIcHdj5lxnpslB/T820KWUGm7IiLbxP7OOhxH
PyUBDHULg65lHexk9UtL8Yvf07jgOA5q11Pxqyn/ofIzbVjIi+waS9HBV+8C1872k7qE13NeoPI7
VRnHPkAqsYNIyW9Tk7LJFu0XXdnENimGgcJ0K1/hiZWTXIVjEZ7xJcC1OH9rXlc25xNClNy/MpIr
pEIJKl4ahpJk7W0boZRvJifFx1rRfhHBGt+zEEAVRhUkxY5pQdGYUHDIF0aQLzta6r1ygbMZfwHQ
Un/sFlrwR2WQB1iFXfUjQYqoAt9EOivx6BAgi80xwTE/VzKfG0/P5qUkA4jhkQVIsq4T1Uc0tv99
i1/64o6qqBx1/S0gClXYM6o+X5pFrviAMlCrsWFPlJ6HFK2fD5h1XbcNc02T0XM2ODrtqqgMJqed
VMp7N4rsWSzUaFBPW3f3pqLs8fJdba2nl32q98XnN9WABZOfAaabpscFV0NsOpCYkciPKca1381Y
6M2eJepZRROkLe3Xd0uUNXVRbJZA/Ke04iIX+IDS6yDoMyQJSb4hKv1uOCIML7RpINKKl3/mCHyi
gXUMK7D3OqOskpe6lejYZeyBb6YoAC5gH15Z+1qV5yIFebirLib/9mFwAfWXaTyCRq/BKbt7UjsA
rKHcn3hZY0hGChUhuj5RyFVt1KVLERtJW8pS0/YjFyVF7Er2CjBUojbdr+H//gMb/UoGA72df7KR
T3kQhpv1e+qHsIjDNlNFErMRJOGqEL7gb2b043/R7PUmDnMKXXLYrAmv/Q8BjCYybVZaN/vGTZ8w
rraA9aeUb0cSltm8eXw3HMRYG01eaArBXrFDjTzlwuZLvlh2KOimpfwbh5Qxm2n719GXY+S3qz3/
R72FYcAZZlMVIEso3+oB3y/Ohoy5e69z3LQSAtSGQOPJ8TPEZHRgbf2kFBqa2FdkkI/SRXgE1iXR
JOCbRM+qb9yk5Zh57693Wf7rXsfav7MgRdgFUwMpSfJcsjm0F65bSgJq9B2N7bjuWpec7xWRVm5N
/uKJCT3HceQt4PIxXXfqb/6SX4aZCgrQoQLF37j8DkHdYAxLnYxwqH4gG6Sf/DxvA7DgLyjeO++p
J1QzMuUvSv/Acu7xNpjSRu3AGVPgbFTM31W84h3mMMS2g/FEnWDS4lYlPz8mvbqVOa0ZWgpvHnE7
yK74KCVYUJvR/wtPlIZ0HjObGc2ieqz8VXMPT1hrVw4QEzfjXfqoMr1CPeNW4c+4TYc5vSsNoxoO
2dnwSSGsSfU0RcTgNN0qvBEWHh/9Zn/SB0OpPcPim3HwpdlBZDTlYXR/nFoad/MJmTVHhp82oxk7
V6tPLU/nXfw5U8yxU9hu8mCgdvfQNsai16lhSALYXkc00yuU/SWDAJoZkoZpTjgc9Yz7m5+iRPpW
ZsWMwd8nFx+/x/Cu1PX1hpC2ODdl0YvS4hOSHmkkwwU/OoyMHeBWDG1kTuZ6nDNt0M34ZX4bB2i4
G+1J00Kh7CQHPWgmT8/Ng/HXRcl+V3sUZCLaiqCXDXQ2t0gj9Oqqf0sOCxsIyuKKyx0zeHCQMRJM
Ao2AqqXvJoihIU/vPVZuD2AB6C7c/9SpLus0zq4nimt0dLYaUyR/vFG4Q0snYGcgR75xoipY0ak2
3nLaz+bErFGHX04BKKLNAWdvUmafrVvIMdqlvh3cippOhjrEKtaKFshSBa5xJnPnilcLL+90mUrI
vC2TisseTZhZaBcD6rTqBC0+pZe+R36mx+beGN0Rz5ziFXvA2zu0naY34wv06lCUAu8+YS98JJqh
9qk69O4+YzYHRr+GRhj/0Rcm1HAUI/Xi5prmslcjwfBXTumq4RtvtVWVF66d4I39hRSsDXGIulxe
FKvT9v9/SZ75ddUpxkaJ84RaCCSPXhSDKLfMhUj34N8GfsPx1z6jnXjl3mVGeANouIuA9iqr1hDE
L5nqvHI+cOyBDrBARFCxO/D3fy6F0fXsNG6nwch9UrUJwycRwVwTcnlXr+5jwpVdNR63x96h8r0h
5sOI40Jj/RKK5HecPJdwKXfZboHqmBmeqEoldnYzwxoYbIV92VsKyl0Fm1FmU/O1egIHCvp17NJZ
WeFo3OWQhoUrvn1Ih9Wk7N60nEC/3toxo0RZKAXMrTJ9RbX401PGKauojzcFvqPmtRXAnHNM1oeF
KnWVk76qbZ+TZj+ch2NTp5WctNqMjqg15t2OPOpkRfpkala/aBPJsUg8qmHcAeV76NSWSaJ1Y/Ej
z0MOHqGQuasPD6bKHdxttL4USwRxxMd63aVMy47Vd7IFfECX8nlyaUyW3/sBomPTvdC3E2Nb3PFx
FJSPzAh6PNaSqLvayd3QXhrSsgcXW5oeCOF3ejy3Wc2op/ccs+bc9DW9xIjARwHdwiAmhG2nPoby
PWHaEo1ziGEcZxZpBv/lHME4EvYZNemMoFzOyuf4VHZmcHORMMkQXIgASTBiPNfHNCwvqYMS9P1J
PUl02bKbRpf50p001HgJ0/C55k8ynxLYJ6INgtGFkqmf8UxCynYui3vMl9pdL3bGmf+Ja9X0ik39
zkyOD6GQapmsdBjpz/A2UQ5svZrq6qYKnoacDCxnsLM7TAa7APwYkat8p8T/fm2scRmk7Uzafbs1
N1/tQxsER3LiQiJFz3P5euBGkozp06/Hyll59UMXzrMNHEUN4wmxfTO1YyDnvcjoDlwOMlOuhW7y
Or3gUtGVlt8qlVQtZRA2FWPRdupR2/u8bT+nNaDvmaEoykY0C9b7QVnU+OklQiIOHk0KrqlbYx2F
1ogDHIYa4PdmYPsDvvHUqsFU3Ojhdx8OlASry7NP4Mgzp88GH607MiKhOeHuCHyis9hnaGVkUgKk
32KLw7DmH8zJRHmYuXOFTID/bu1RCMLKAGEe1hUTXUzAfsUxoc6h/DAh9hSZsSXPdpCJIO1XDJ+I
31JFxn04eoAj+tUYYr/HOcdk0ScdepGKUeTJpwUbRJRxFqeq5jWMAQ1lDVGelo7ddDNpmR8pSUH1
oNrT9hPtHMnFDeJ9gOWZvm4sIgyA9gyBY+8bx3GDZabTubsKTXaS8NRuc2aKOBnbCNSHXnoo/o1j
yfTntDZam0FeyAh45dJhBJ177AFJ8KzoHWXnAtZFJOpf86wMTXj7nbabHfr5wSddoE23l2a5z/8u
RjZkVwi6Z0u8Rt1DfmuJ9hMJvOO/7JqzQQxMrTJdr9TVCJIMEqeu6G1QgDPwGnvqtw7golEXHyrv
HVStuH7x1epl9LMStVxn1W4STyLiU4XrtP1pMc4ivgI3mJnKhbNTPQ8fccdEc1AkriJvRLtwjlES
tv4f82WiuIRzepxw5eAbq67aRXrkuYtB9B8U2a93DsfYPWTc9gJa7JVxAtlN9rYiMtclzD4hQ1oR
zOflveqa/9YXGpg+n5KJs4PRgwHKbrvjyprBcGOdP84+3exmuTV0ttJhhL9i0AyiiUvgKZx2lAQ4
1bMUv5XrZYnZNGTh/3AXzZjn3M0oKNuQFSzhCezMKs7930XeUvqP7E7IPoxINj9nlS+vhnedZEY1
xcN5yVAIfd3QBAj0H1CoIgYpe9BUB4DfSxtxsPO+jSojrpMySMJANWG4NuQFwkb9KuA0b16mZ3Jn
NuQkRV2tq+eD6a6cJPUdMOyKqA9mXexH3LTfEtsiKXKleG7yG3l+ukO4G3z7O1ErovjdyZ5kbdKr
tPlRt2zyTh7HQ2lMRI47P093PI2CzjNjz26wNl1sCPoJwD/e17pzf+mFmBGOpHoJM9micZvZ+4Zc
LlsBZpE3MLKWEy9XAslGzfMT+BbeksmIAcdU8negbnaS3lsx5+7RZFxwvk5ASjcOZTCeFZYWi3A1
hKIwbJyPe16RddsIk28cGSoJ9zUFUWZuVjLTtcNa63I4g4F+LovGJe4tsnq1EEvods8e9tdu+wex
0QBBsCtCQ5hSrKpDJ6d5tliunblz2xX3W2kEVhUCj4CGiROQjPJS5xquDm9yW52Fndy8n6vafTEg
kRmP+OvAHzVAWTFHS9as+hdrKPgMkUxb4I33pOzR0jQWMLb4ayVWkrj7NMogjpz9zLmbF6vcTPfr
6QkY6W2uAPbaYja+S+2OyaoavWkLmXyhbA8+89uABmfCNdaK/39VYJ6lFU1XjWR7MfA+cSJJpTPJ
xna14RL2AMbj4vlLvtx2DLrFzJvkCcKkRyvcStLNA3hT8f1w0/H9KKHjmQRmg+fwHs7RdG0e/wdT
WYLTdODsaO1UACcfhXggd60Ip4zsvLC10WtxdCByN5QtxX0p9lTNiLKBdj1DFRu+JDL/hOQyW2cn
Y5GXNhHQluPqmp7mV4FjRa3hNRJCX9H2dG9PxRWfVECZvz7G2Yx0oQFH26E/7vZTY0bSNSUAYJey
UiCjtS+32pQF4USGQmN7VO2ZzEDTWv2cyktfS4mIZXmm5xvdBn245blMEMJPCJPTHPJn763lFVyA
eqZ5w+z74tvlz48xoTuqGsA5jNCAqOeCJc3FVcsRB6JkWFDyA0GFYuaz2O75AIPqcshkFuSrJyz/
eo/dJZ677+P+oDX11eWaGcj4VQ6DP05V7y060qHkB2/zJXxm+gu/qsDQTalA4v/9UKtF3i3QXFhy
iXblUhBfz7vqs4Zf39T7cbfVhk75saU9uYTnmJrrdG5L2l0kKlaCuJ5r2fZHcd/wznCRlU0O234r
haeq5vXemFB3esLNn1DCsS0j6kZDsdOTYD4uw2iTwOsryFivns7ePNCaKRoxOOwrwL//ZqxCK3O7
YM3v7cZuxFOgh9O0Q8XLUgJ2BQYmuJ1256KYgmuGMfqKDCOsQSkRozH7mLPEBKmTQLByZ8WLjo6w
C2wrUL9lQedj+xfBEFJIJT9TF4UT7QkaZfOzay9H/KUPd3qgID6ZY5aKHBtfUIlGoPYp2D0ULQKp
+He/LpkNhzgQuLAUYjzPBtR0uqmpHdJsUQ0l85luuI+rZa1A8YBTEOBMESwlt93KlPRvIFakRPCE
dmLkuJQnd+JC+p0spWEzBdxWooP7UJ8vZFMtTzkE0kLgRqNoeMkAg/ZthYvpR7C5mllVFnia4SvQ
yW5i0dbUorXci9nrzzo=
`protect end_protected
