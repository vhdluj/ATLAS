`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kAXwT7d658QC1dsfnH1QF4NIAoz5+alkSYHBTRtmerS7p1ac1AO3NO9sGPgtlGG5Aml+YvkMakZF
/szY5YJ+9w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ozzvVs5dmDk8CJpQpBpAcwD99J/dT9rsyFsBlnF9aRoScUinm6CswJzpbfwfu0mbfLpRSJCke+J5
qf7zw6uMxl5i/xiEwEW/323W3blSb7pRNKfccRxFdWK0XhUqGOQpKwOqhOHA34u90OyH8liFaiPK
nPTR2FRf2zMncpDE6Fk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I7EgujdEmHQlV9LUFNPZNiBtedxY4eQjCs5eA3XHObzOnOW1nfLd43osE3wuHXF87CZVIT13s3et
gdb1FbRA7+8R/SzYYqeI+VHz/HBq1bTVDxm8lD62HZLCoKmyXD99sb9K7MkNpOyGF5LzofArZlVL
awRCC0tx0NKQqRTE4adedFgTJbrcXmqRBpzNrEDE8jn9fUpgk96L6rFoJup2WR71zr4Y4NG2LRXL
dbHCDOEwLsOMtDq7ItrlsArmhVJ/QZYTGPbMHiJ83sruG0VjET2/betTZQwCwjGhziLhFr04etRi
ADaaJGbyTyqQejTT1GbKGQzVUwIMOehyYqVJVg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NbBpnMI0YS9SKrPVaqHY7tqNP9e6ok6/Y4FXS7GhJCM3zPfWay+W3hmtw90ws6BxJqYHOBf3/Obw
wQ4f38fIOYRfgcRLTDifgExsrRv3MLMmx2Z6zxorMcU6vwDYXE3ZW+FuMeiKM8jdvtNLAFKlyIHq
RXrttzAwHbn27rROgeM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aZVl359rOZyi+ehoO+iIlq96VOmtxobLVHRWdfkB9CHWUByF/ykacD8J7jzK1AGHONkeL4KYsqt9
FFUnZ/yZTdECpo2iVTVlEz2zz3GUv6dFtk8FE05oQ0YlD8JSA2+MBqCn1Ts9SMMG6T+qvb/MC/nx
HlNBhtv6nzdesmeXvVxYlJuQWLacrBd5bCXHxQKQA0DvBMFnNY6tzXX/bT+hKgWPlmtG5wUk4EQI
uJsoh/HRKeWn2KPf3rTNy+Lt8iHlCBxKl+FjdeRckDgSmqXzfgywbFk0CBeW5r/t/gadfvfnlKTu
wYpq2CbDGgr6buQcIqkDrNxGzjDaYKbQtzaWKg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20576)
`protect data_block
pAJy+4hOtBsWsRtEwfSJbJpUm8443rBj/9B1dcTq2o8NCJzwoXTTbU0OBSmW9nmPvIbVNFYvYzsf
fqiQAekdpf1RcsyJ+0DiykEsDHV6Evj2fuqXH8T78DS8ZJgEYBVpkwiQBUYeOP1O+CRx7uGhI8Cv
qWm3RXWiv1Pul7KWa9P8QVX6bNsbvxUXlPZ+KlVyH7I4DqYg4GitI6hkomLpHS6s+VMEyshQPMe+
TsJkJnx13WhvauQFHm+s8Gn4QyYQJLufs9lt3TK+gNDF0oynRIBfEGk/HOvfXacuzZ3dtBIYLjJZ
FoQAuCeJGXrqkL8FX9lr0D/0koyMHP35q3K22c4xcA5ws/xbH0NmYG+GuIdqxJcIOIR9/RctecfO
ba2LneTahaikEdvzewY9SEBxCPRQlEV+0fgeRLkTE3aIckbS9wOy74HBPWOyk0ME4lwV3KsdV9oT
81Ahp2IUXphS2iH0ln+jQzmWAvLeOEuIBGriBFaWAR/LY3jstYogiSy4vab0lQa2WlhOtuyLLtRt
yO3F/DRX2sCVr2YG+RpsFqINmvvzmBUjHZmqnSYKEReiEp67EZpLOhYVhmlbIsZQQwX3v8Hn289K
qoKP98OCkOUvwxGPvQFI1BN5MqWAgSV4poKoKBr7W8/2xJQm6qaoby2l2sLpln2IRzFTfkJ61cvn
i68VQJrKBRDGqkDch24QEj2eiq3C4UzYhiLfjoNk2BRVjPGITU4aBJCNko7zL2EOai6AClvsh45A
WBa7E81ugpxsQflb/eYeg76x5TT6lJPuSDgCobnwc5JBBCVviPF+Jkzfl7WdcWdKE18IiFjcGoVp
b34Htwfy6KHUSWvDXzxheuKY5hCUSt9DnIlj85K3c94Gz/PtWblgQ7l/mv4Qxqwk2cQLCxIrrAId
iMazf4vYPCdllXJvLKv0bqqbB+5qtgvMNKxWsPXi8omDYyFvU6uYQUH33WMbaCVRcgU6uIOL5G6O
BxXNcL5gq+Ir4GX3sgtR9cRr/lYXLD+7pR9lB+sbIblhiraBS0z0XRpri1PWDMaCmORFDxBEMBbC
MoKpu3ZD8GheKsacOJF09ZhdDtnxu4iVZEEclgOjezinqNH3jPNls1Nf0tKG9em8xaD0ksM0UQds
RF8wZHJ4WmVLYwyEN0emOmsE2ACHSxDvF8491NmV40sqHnnO69c6AQmf8E6zcIa5pNxdiO+nQlYH
S1sxttoWkG7vrA8LmF6nWhN6iFK8Ftg7I1LOS+mFNv/ts986nKNoyDuSmuvSCgqeD1OHkIlaFgfy
39Zd0zHiHSLmPQcxL2qBl2z7FTg6X6Kha1lwaGhgkXgX6X2HD/dYf+dzPFNLL2SJe73MLlfu4/5q
TbR3gd1UJ49Z7coFUz94yvFl3Q5jikbBF7pCADLro6du3IvRw6regxX054lWTQTVXlP2ugmxyvB8
09qTSet/VlsN9xN2MnSpMw/kymJRrpXGZ2ocf9dtD+SGjXDsELlgdemCynIO+S0g5tL/wcS9OQWw
nvIZRkqsRr0s4/pmGemJrSbHy7o2/NZ9ovW77qnjieHUwGwSImiwBz9iznfEBGLlRHjdjBKDkbJS
XRKD8913Fc8ziiCn/NP6Ggj82pgcEgCNKvlPtDpgxthYvbwNOMSKWqpgkEsJzJKnxj1w0zaForhI
7N/Auiey0yH2EKc2XJn/YCOi5awGAzk7QOqKtYwOmH+e4dlcZegsK5eVOIRPs1gOIBXI8CyxiJxk
AjzCxkax9zv5is/Vo4860SeKZOOO6NVZ8sqqcIsGg5vfKr3ApkvQ8dImorGyGd05nfPs24JnQ9k1
jaYEHUVRbypFi6qrfuBczzUkf6lNFpoy4OWj5DCWgksarbTv4G6S4Y+Y+BueWQiQdFB+YHdLSDG6
TGuYIguFJ79XhS9OPiEFtHj6umiNGl8JXdJq8WT6yGPVzRVwlS1Qa89UhXAIU6blKR5nUbiXd1ne
d8qJvFO9O8nByPYJVQvqpxz79UZdqlyILrkbEGGW9aSnlul8tNvN4aUyU1FxG2kj+TFmbhLq4fXI
XxWS3Lv+yhnjtBhPKzrao98lj8t+vk0idmCC2B1CYtFhKoj5XJgxmbhNGTygr78eedR3Hb/2N6hg
AY5Kz3hDXCeKwhhhJAxYFyF/M5rEazpbH26BiErjOpjNmOirTRK5KFG2edWgAgBT8jqTsb6Xsvos
6Irn4qbjg+0j9tYs27JiBEvOkwJukNCow4JS7q7O7ne/4ePsUKVifgVdB5Ira+sDvd0sPtyBhF+Y
bqO9Ds+rs2+C7FgvHCr95POAH5hGo4GDW08Yr77HlbznhQNYSMT7mnss7lBt40Q5am5oEw8pP+LC
+uyEE745BJipWpk6Fp8I9lzd9ZeTGoTHyqR7JqpQ/H1sXhnUCAhyymTv0UlPzkBuR7P3eil96IU1
R+DoeMAi5Cjo8tITQaOK0QbY6bCp6qn1103Edf6sGIldyfIqaN1dVRDid788/Z5OH9JskGWYZN9y
60zdeSwrKuRV5SGBlTJ5YiaaXwugQM6wga14CwX59flx9D1Q6hZ/PtO7cLd4qIS1tjLvHHiQFYEK
xCWWZdSP1ohLxV1ZydchIP6JH9hDWoZYIrSCoHVPzZCzrH5khgWMTrjazwEXrmaapaw6AXO1kAE7
ZFlLLZqX1oPlAVgldnFUK8Ra2k+WWA+v6LwfUrAhBAp6yFvG+69bt3ixV3dY8ZyzCiCxR4Sfvt5H
0Xl2tJZOVFpVT93gO0nx8SQ6Ya1d0u4x0u8oOXVrGC1r7JqkxDrUAiaYp3bySTZK8nOkrYbkhrI5
t+qdA781MZixO5uQQn+7LuWSpq0+pIMKg9n5F3/gDOwYdhMplNJSpECSSnwyDjxQzFUPqLrai1Wo
zS05y0LCQaYeSR4BSNlomCTNf9Qx1FdhirfuTZdB35lgONsrBmwGAqxVdYhDMyGL2XvTtJJP/0dG
pVIzuJop7OJIgGFJWvMdAeK7seURAgJ/7pujnvC5g2+cJgX5KVlPsPJOHLPGbmy4Cv6c5VZ5ygXu
yA8z2V2SM5HL2uyp7hN1aBgFwShzYTesbIElWgHi6AF9ofabK0sPFkEz7cnB+zirLNS2/YT3jSjR
XPw0ybAfejfl4smE6s97BGPj64cloJkzhbhPJM6/ddg5NjhEOaqm3ARDB1UJTxtL0876FJmGFA4u
iDauXdH6DwgPUyPFJNd6Hnfg5OZYyj8loG5LzjMJi3dVEg1rPvW0mtQCxw0JlRX4Bvb9Kvh9zzVw
WLLK0fcYtwvTX1l4NrQ6ND9nvro8jqHhax7HwvRM2gkfeR6KWYJdSC50c4CbMSWyZ1/JeWiSL56J
NJkZAOESV/NLK9wpGbudY2K+Y8vdRE/62TqqUTcP9OLmVtvTM7ZqhXf2IeVVtNNORssXSk+r73Is
I/0NHaLnOMflU5vFl5Ae4P/loOu4QbQIMMyQJ1ByLMBj7Z6+X3O1aP7k4fU/cegatAEgc3FZ1Gfy
lNkWzX5CII4JXdvek8LHBG9nk/fVmXrwQkBJ1P5SPAmFIwDt5ON/soBlmHysYuF6Nqd08GYF3S/d
hQqzIX9F0jgENbIQkQMpPt7i/E/0ItgxB4yHv9b0kJ+r9vwmD4UV2sBxBA2HvJueZ+YtZip0vv/c
SCoUOemjRRpjVQm9vKf1bjuZaJbndYMifQxjMA1p2ql6b5nR85MQpDIuRx8Ywu2pVR48IkLsJlxR
rtq2ElPukx06hXKhpvPyJEesG3l9me/rH2D9JP6c7bEeJeqUSjoi/RknRcdQEozWnUTOdWabthZL
wEmmo3kJli5Q32izvJUii/y//wGS3pIrdjf91S2dnTOIOzf5IRsjtb0b+tlONW2NPVDHzUEuCXjP
XrCGRHCafRIhZKyUuy9qlWcQPrf6yOn4C2p2FMB7Tz93EXbXopRlNTnFfC4RjjmnNjNDmYM+wesD
F3LtjseLym62uOwLEsD0YrLZlCHWTDoYb88SWb1c2nf1qIRReRCyjMQFE7OB6VEqYfp7Pufl18Xi
B3raTDVMxbRQ39P3B40dIxTu5UOeMb9iZTj3jRwOrrIOb4g5Hn1I9/G2oAef+VwXz9O3u16ERvjT
zsxezmPzc7jYUSUBe5rmYRt7JhZH4orLITDaxGmDrN2Ej83j6xUlr2y8gVtueXtXHOzmX7hPvH1Z
/GEXRL2WsW684CxDb9Ke87L6fo0XOp0Yb5lpbMA/r6DBL7by8h9o12dVMcSrPHmK7vg8E0G+yhSh
yIEobyz4DJ42zk6Vx0fcZXRUz2Y8brzHUi4ra50ECfBQn6ykdGzD/kRSvTAp9n2xVdjmyGAB2BfU
83z6L88XUNsVnBN7GdW3iwHmLCqTaLdMoQbmgMLJFn307ArZ2f/OBJmikdKcMitxyPuWszFPbABb
ECWbson9PASPFlAagHa4zDfHMRYHLtv+6HrhpJiTDOVItXgauyHc57xcEYbffqdOgZJrCgceq1Uc
WUjYdA7FvZBgLtQquP2mR59FcErosvqkzw7jIDYg9z8jPMdBAOwKabwOhlt0BzYl2K+h4JDfLBVq
QIBrxZs3NeeVLNZrpTrbdiS+UwgplW7fnNSeMvf1tszuwD1oCA3Delo3j4He4L2F8B/damJ9Ua9K
kHhiYQnr15/Cv2IfjLvYYunLR2Zt///qDmPb7nRGuyLmHD66OT54AtcsRzPLYmQAE0UzmylLm+XE
bYxW6mIwbdHJBBOX7u4FDOoVR0nTNX7a0bCuzmtZ7GnVyopQs/r0mz1awymO9iZWnGlxeOC/5HIG
4pIdy6SnRFGbXIAX2+AaycN6jTbPnMjm+8znaEeRaIINUUjyNZ1UIVbTOkuKuxIyLx+lvO7uLUhe
vLE7YT4T2d4Z8aR7cJz+8bVgh+nImiqtsKL3nWb0lgLj3ox61C/9zVr/AbcGWbFyiBbqlCFRenWS
JnD2ZbKFZZUBxtLC6/WSG/namJTliYLJrotjF81BkPRctXISICx2rIca8ymh429FC00kSZFGBRzp
OdFGHlVxWIYITWjYuMYTzrO1hmdOYJsgiPlgUL85hOBNp4fQpkY+5ygiLQsIj8S+VYU57SYoOrw6
J08eGox76XbcryUGHVsJtOfznab2sk52L8SCAMzNv4SnPv4eu5wkkowvlVl/z5IMDic1ABIri4Te
iCLCv/I4Wvkdm4VgcWHMuZ5l8zL/OWodrHXwaQ2AJRmjn9VjOdKBDGv2C96tc8C7id0vy1tV3/39
u2qNRd1pi1rQBhR5vhkbYmutZP96F9yUzn9gnRDBl+EbYCdTLpoMiB3sLTl9m84nFLbx9yjzCUXH
aZqGD3tLO+l1n7y03pWj949PnrMTPH/FED4J9g+KyMDHioSkKe5XyHb6EKucLLIbkOZoVNk3Hjy/
aHBBMRPzIgSYlTCvpdgZW36iwX4fOD3omwPp5QId22CH7lv0+pOxak3kF6VAzOpqzycaZsx4NgLf
rGeMcbORmnZJYOlHAxuyRLnw4dmxnhNYRIuIaFOC9y9r2V6oLkKVCt8+z8SJBlimhOUQrHgvd4Nz
ZRditUSlhjcAnpZF4fPp8tWDe8Ssqij9G2fO0mIhO7xB7KzknHW6Mvy/1YCMcoRYhwlD7aFhElf5
NIZNE70VRS8yeiIf9G45Pvg8irOBLA0vENW3zOXw1OycEDRmx/PTV+g5qsB0Rw/PvW6G/mOWrfHS
2TAcLhfWyyjuTh+Ymr/P+MG3t1qd8aIlCnawvhQ6CpHVgwnD5iURJ1qw5hQrxEJ9T/ccniEIqyBk
sMCsIYxJ+pa2X9BpDJ9TTV7l+12+/CrCtpvr3awFKBhd1d5LYYsMcnSCRUEECdMq+r7adLE1lhww
UpMQS/TjteABmrZeu6UTO/8JcQYMuhQmeyBrgrxu5XekLlg1RebhTWHvuXDN7jDcrj7AUK84sm9Z
8Cu+RTXWq1yLs1hQnjNVFxZag6+jxonSehIW9fda6Q0KZ/KHUV3NYdh0xwaL0fB6UcIuZbYvI2zQ
xxuHa7i+XfT1SywxkycGGmyFxLBAD8xn33xDxiCpxby9r5CaYNnBRp3mY29VsWa2ILf5MzLWC/pF
a1cSKGUCyFeFk6FRWKciF1DRFxUmqYQhTuP0QdajvRUbjIqWXOrqBfUjX6NfHsGAjSbLj+cLhrEu
gNPoQQSrqmevLjnLT6/NLdmSU9zb1QtAUwi+1SJv2w4Phn0rROF3PbxDMYVkKwFKJ/5njrbhyKsP
oPaJsIUVsNAftelht+BK8kiUMVJfiaDDs6TfZUfHYy3LRE8184I3oimtLwJrsN74Q8PPVfK6pS2W
wAveHjxqXAjjnFugLMFew0Hz60sVJ/wa2q7p1AinKCFdXAp6dVnkKNu/8+LMWIt3LdhZ3V8CkPtx
tq66c/7t36iiUQlroVhPQaTu7nc25vPW9tkzqNrSdXTC7LCTaqqDZKugJ3EZm9qnc5oQMZG6FC5a
BLO5+cmBAjYmtbqa22NKmNM7uEVR+44FQ8RanfCbAFA4HrU3xQwu8XOymLztnwfSM9qbCRPEcF9y
MnBk4ciAHoSy4H7H75MVTj0+MXGqRgrYion116JXwh3NYsFL4aekEannR0mE7dR3AP7/49FWZtue
rxBxUHPv+PrrGzkf8YDQH85mByLfwYjXbgyV9GaOoPBuqv9CsypfvEe5HzHla4hyLAz5O8UvbCnJ
FFA8OphMyzLJjtQLSD1OnyImh/OMJGP8lDwqgyPLIigJGTVztQiz9t3LaNZt3tde6LB4ViwLuSYa
m3TqNbw56G4PH7NVVbzJju8eIDIhSMI2wDWMoHa8K01jcyhF3kICG5d+aNLq+oSg44m1ShzNbWeE
efgMoEjkNYt3qGeD35OWmpu4UjnuJCWORa118B3oJoDOkDznY58Br80ozLbVntj4nerYUkEq7Gha
ZrQiwk//PNk8lN/BrqeLrNH1uWmS+A9l+b9iP9Lx2zv6ERc+XUY0083io2kxe112nW7dTz5RwDmB
0aeRphXKiwaIn2OQuy+gjT/p0Wkzoq5R0K8mbnRZTFk9VQSZS4jONaZwvZyIAn7USas2UdEsaSTs
Ag2Wmlg9X6NjOkBGxrsflvn+Q7XX1otvvK9eCq4d8TwzVKHKfSXjWZObcgsE36bhNbVrLk18I5av
5VFHzQxycbXqWmfVwlXEZviS9j7tZkdWeLPk7o570EZgdB4ZzfWVQ2bU/A7/6v/9QnCxYZpznLNn
+Bsgs24+pE3U7clgFglRKSTTusnEZfq10aeXWLIOixMoVYPwTE4ymMQHoLv6dfvuBMc9TJCJluVJ
xrwBPVLU5LUgBAsBrPf2ECSG7hwjuIaY5NKGg7ZlIOm6Np0miR///CTJ2qXBwDvpGqAt9hA4BNYc
b49q7JpN1cPkWx9bEvCAbGgFngxBFZ5m06eZ0V2IiCeqzCMEzmPQ/q2dYIBkOEC8ze/utBkxWjlg
x4Y7uKCH6AALv+blE5bmYk/XP8gF/+9ZhuKrzijJScwQK+mjfeMESJ5CYAsSb9WwGTKTAiE93iII
VXELwh7sWl937qpiXMiwHYvhc3EE93DbqhiPlbJyvK4qn96np5snKDECVNHlKtpFc0DuUKBFo4Bu
jfy8YQ73K2gLfufGeevavtD2bbI6TzLygfoZadxN4lPLiLTBjvd+eesH7OrZZ9UVQ10SqaM/wPg3
5TrPZsDbuFs1ApOIA58MlU9/PqkpcsgtdUnbw/vUfsCCiGm0uud6YebDKp/t07sdlq1kUeAxtrKP
efQsvI1O+uRNe4K6ghtWUrkrU9M1w3Xza6/9HYr//moFlbR0b6TLjmn1CFB3nAEdP7H1qzF1Qyvy
hMye0ekO56089eh4aO8EKWQ3TKqJSOL3K1Jae7+jiT8Yn22qR7UV/Ngp0HkyE2Ausc6ZxiWkWZGc
jS/3XGPnGjcBK5P+rdUNaSXapiXiOecwSmOBWqH0dLyJ9KZT+RgSYc+mrUXw+pF9/sCM1iR2/0Q5
a2r+WVUnNjm/O5hNdW+I4w3jmBSbQcefPD+PL86kGKsetpludeMprPo9wNCRUCX1+uhNLjICBo/n
i8VzAYckizjh14EHhOpj3+43mBPtHCZr6RadeijdrTrRg907AkgyzxVJWN7rCu+6MADw5644axGY
rMHBbDIbT1mS0ALdHfgv+gPuDz7aqLZhnAZIeFQ/67XroP1KfOMMdw1PJQxIioKBjJEWnghQi1c1
95mATsuPnxSI9i7iW5aBZEXUUoCWBx4lJVuyos3OUXjK7War3zQvwszKPoc3kkIMFCnaFPaAEJ9N
HQHJdHpM3oKPM4cSEbMhCduII8wvZ5tQCdh3wPL2nSx7yFL7roGoOP5a8xdLSy96nikMjGxE0e2Y
5gDOBGy7bytyqpmgrr7kGAVHlouBuztz7IZaeejaFQi++QRWV42dOGnV59a+I2M9dsZ8rCEnd23M
Ufueqy5eo+pkjeh1HL/UdAAWxkSbRhmcWKyVsUQ+fgg8URHcTIEZWqELJpVbVVGhjVan58EdC6AO
2gRDcFvWIaghIJ4KwDnYQUoNHZU15Xy+zNAojXRYr8V9wnaF3bFMtIfryYcR4vWi1YvU6ViPeTZe
ClGQjdonkKm5QdEi185Ni0NnQ/cjNGH5iMdI8/+w7BPrBT5WPLpnFpoP53lNO22QxeL8ARBcDV1E
qAcATXvvYrSNQXOFQ7S5iBytPmzHhxmsyuBN+4iYBlsNumThDs8T5SGUHMd7EmgS9NnA3csKy8c9
Z8v0HJbCiTKdNL8As59sO9hnqRiV9ykX92XXyDMaOTjXNLKghrWAmqkirF9XBRMTsdNfdlsjUPZd
kw31/VFo6GwAyqr0bgY0258ha+WftwRedhakDH+yez2VKEClleh3P+lHy3loDgDBYP1xMMzoVcZh
B0bKhvahi/+klnhBlWSuaho+H+6Pk4KF8vs2hSmanX9Vgi9BqsiG4Uz5paXPmCzB1wBELtZV96Dk
o/riondKo+HBaoYd3gS6KL79jNH3GgH7ogsMh+gRed+j1Oiyxwuq0NBsefbSOpTVYnFq2E92D5I/
Clr9OdPuhTbRUGxrWKhCm7jREELWxEQHvzJDazizxa5WwqpX9skXXvqaMje1yTR6LcoRLC7W6Udl
L6dptpQFx9pTTMAgy/PFlalNMH2kjDOM8J74SqF0TDhLqfouUFV2PLwpm9Ph9jzHUeFFnpG92ekK
JwFPqCFsCMMXYmigz35CmTdyL/LNBkAXHJPV2jhxy59hh3/o18cI/ahzKcZ/f3b6lGIr1VeRJ7pp
7nWp4/9c67Wx6M/07/wcDS21cZgxmhag0XfQA78UD+Sbj88OQ9KQuQ1RTcpkrJw9DQAsvgHy+Bad
lOgQK9Z2XksGbH8NFaXVpBZ+b54GOju3WjNbGD/FLKYLuK2YnJoiMPluOophRC2/H3KLJmKhmjhn
HZQIkV48JNoCJ6O3m5R5XHTefzoAsBxsKI3ciMsUzJBF/JcVSO5IouRbkg5lO6C9QMuLAG1BSe3q
61TvGDxm2KV6C9QZUPXfu9YGh36ij2/Xl+TVL2c9ptxxyQTVDmkW9rUGBF/ib0E2o+G3CpDlalO9
RFmiEAA2fvSszebsGr1dt8qqEcRitvIMY/cvpupgZDZBVc/P2hkMnGgxC4G8ll/2fod7VZ2A9qa7
6L5CLm1RxKoYIWtbB9/U6RPNsBsG4k86opV/Yx5NiVFOhsCAZvKe77RZEuCdEwJKweCT89DwLDJ9
vNalMSsy1AAMrZ/L4RMCpAweZJCYhIPZNhSuC25y+N+li/lqHan8oMKBYhNqNJBfyAb+foq6OfBs
gZ6zd4k1UbUCcnETmoVpqZaWeuk19gQmdYyAWI248FztvCpbytwzyHY7cHQMX9qU5TTfplAcQ5fR
kpL0lpOQPI1bY3JeuvE0fjif/hY/VNV7KxrjiRAEMzAoOqMOk2vAYmQfgjsSkWchXD7183PvyDzH
goM11WEnJ7VNuOefX4DTPLTbIOZe8lj8kv6iFqfLkanmne2cVMWGmkUZqGsA2aaZ2Wxfcrj/L5yw
os31IWWNK5TEjmwv6IoZSpBdSw8rqn5K1llymPIEUyQvUbRSTqh+UiCvShPQZCGjCNSBDlQAy5kG
xdvt9voGf5tb7Uvp7Rqn9TNrhxAjvOhF+n8R5WAimgksMGzl231efpfTbaJ73pyIb65h/ZECQvbE
eFhf2kzNmNm11WskL32QErZYXA6xKDR0R6l2HDchjTN3qn9bCzQgQ18YnzDVYZbkw/uk4sbjBSH4
Az/8BO8EEqEBP11jY4dEYxlmJh02oQqzj7iWIAWs9bkqAm+6bwLqhxuJDc6kstYesuW3bgFmODMZ
fEDqx2xGAytXZdmopPSx3mQu3JfbiokoWCapEaodpLZdHzZIVIwxUaf+5eAdDqUlPqUT5GF8+OMp
lxJgl7eKGLfCz0o8mC1s2+wcNfkDipx0IhCq0CGDsZXb4E1RhenpKscbj3jnHmIGM+XzxOJMy+Ms
5jNFgaUtElEz0xtXO4xzL46zOuNxb6Bta6/7O4inNE1L57VPyL73AgdSkRGVl1huhUAW5s9jstB0
eeJZMe1bOD97Ltcoh6kDu8WUKLBu54VkcStcruEka1xj4kBgK/hR/MJ8UxmNV+gErx9ErQIC+5V1
zUPjvLHuC1K58z+Ygr2y7QxBtA4X0BwV3pRwOeXSKo25O9LZhwfS6UqMgoapq9RUAh7rYtgggkfB
e/wPF/7swDrJFGDALn4eD0Bk+7Hmm2lxx3i0H19mJA8yBGDoFQqBGg/iKHh5o4vcT5wU0BVp53Lm
kyEP9oqCzO4S6pVpHDfIUGd4TE/52e4g0AK9403hy9vVFJ5wAgmTor3x6+LkqqpbgyLO8/4s+eEP
aC6jaDjw4NG5RAuG/L9ui7J3ad335Mr2dud80SlzMX16bNrgI6J2x7NGj/XjkidMFCJ2GEXAKqqD
3jOWeX6736CryzW2ffNQt7pQoX6/27xO+Xc+pEij31dIQtiXRQoTOx+IudAoE5mHguCHbbCh3JoT
w2GiMmn1OwdTUsBXd4YZOWzwSPSE4UqMo3opDGL8Iji69eyhmgzXN6WAf3+BQ543YeaDXfOXBmSK
U+mgeHJlAXXSH8BsnZF3QCpcpUAxoCevYc5zQD69+r8rpwVLLVDeE0F88hN9RzLW0WDbEKl0t6rW
21RyDq649H1N9INhqrBlyuA0YnGW3d55HW3gIMUIFwIB7Q5O+F8NcqlQqM6KXoen3DbVt6vfk4OK
sThv2riIh8Rr18nQBQsm7s1a3TVsnnwUdOBgLOMavWlTnN3hfOonWB5lp6j0a9CZ6Bfq1SIEfFCS
Hkq5L9pxJYqsdNECjwN0pucks4xEXwTQoBefHoxILih3FmUBfFkR4OMzfugile0SQXC7paO9ytoH
xLpE8yIc2i21B3U7lFcbcE67SZnIaC6uJFGPvd7xaj3CgoqVFqqlhUU+dPcj2GYEVGBS0fx+XnIW
jHfnwkNOjR85B2pgpQtek8L1aGUk0mb9NYwuIvfmJGjVU4kl37DFKx4heb9yjpyj12b7RnS1NgQf
7euPe19LGgUPiNohStfLUJ5lEbZ2hLcNajWvuvnK011n2Z5y2qJGMNmpYGwv8N9XLjYWxoMYCf1f
guWRf0m6n4eY4iG02oCXH8yxMbPjNiMExJ/TxdHkgI7kfFIVSUXymQZhuzVqFVFb8ZIsveldseWk
+pmk5TI/wT8g9lxQmE+tNVDEL2e3mQSNHDbU777WSxoL8nukpyKAol7JL/6Tm/869H7EQogVlZj9
I2/bC87RmbcshQXXFXFOHixwH78zdvzdyDA9+p3pQUFHL1jYdDX56kvJ/Dma73UVW7RmzUDwEd2M
xDhlCxDpK4vBypsBR9fWOuS8M7Zi3XIP/3TVUAqFl+MsGyv1rvLsIXWWi918nZM8j1CQoFDvptbm
uN8cKEsKnIUa6qx/7MWjuYy/YSBgkJ6va14zkVyvl1SB357EElEDi6NqGyn27hFqv3yR8esPAL9b
xaNtGWGOaMGB6N8TvDMkh9Vo+bV9Pau76pL3hn1qGou7svxmw1UGiiCM1UpxFMjyLGZlqizGjtAy
U2GbfbZiwSjx58rlJVUXCFHw8rpi/xAi9uhW5JHYETplUJnzYw5bdPogLmLbNlACBR4UAeVKRXhq
y0nEzg6ws55wtil2gfbsZ3bnswZgGYatBwP87jfV7TaLT99fqjneT+9wPUaOx6Q65Ts3SWHfhr3L
9CYdHt+Yovy64rJaJ7dDlubkWKBFd1bK7JU0XYoxPi6MLfSmp+7uhxVpasd+V75L5NTLBiAU0Uvl
TocjlfPzYWlS268ZjFTJ8pDBOSweSaYAHTl340cPB2Xk5+8hr3ERQGhE/YrdtaFwYiazQYoazWyM
iX4KkiuqE+gFc4kLPhyRu4iCHc2vJqVlOQs1/Qr5kG7ccSMvV8U2kidvYZ6AxEqYeniQ0n3kS8m/
STgj1tE/+EqYkzAl6Fbf8rArafoQnkrMcrxzn9r9fMadHIEnKS9a8EjJWQ6sHRuKzS3ZuBYp64/q
OynZ28kVItOZuLWEV6tqd9wFSZlHnojW/HHVHtPaXsKthhfIgrHgADjk4dlYIiecarycW/A+Ps/w
bejZUPx2z6T6TLfNqvhMaYQlDMe4f06TWMju+uQoeF93ADCZHSONziot8duKrQdZci0TpKIgfFr2
ALXqIY0lFJJsdqO+LUc6UDnLaF4p18xMIZBpGUuKLvNQgKSoGyJ0qtBYPEx9zZb2ozqndKWzn/uI
NhlmoTCpVFzoOcimIJpCC5j4QS1kq+Rb7EBPJkkTIn0LzrDCjwrbnIUoI2uEfmyVTq2WcPYMKoOZ
taBkJav6CH/ywKfpF5kmK1HQ0ZwcgPYcAT+VG1HNoHfu9tef9c4LBhjwK3jQOlS7dDyrkDTVmQzC
laUZyePEjBVHOh6vOQHtJAEkWpqBpJ6ycJyF4wJGk2Gp68NgEAnSesbA5XqjBojnL30Va3msINx3
AKgobdM6QzvgSEuB/cjk7Qw/RtGn7pgWRwCCetMj5D7yo2QgrRJT93PqnKorn0RL0G+/2IvYja9r
QAO1tYL5r6LmYliyNxtgd5erx+tsRVX/TQE6dEjQNRw2xpDzbIFdF8fj9B8X7BpQxUSCNsJdNG5z
tlXDxDZ5KRWYatBuNQGR7VawF0LKf9MkxmbQA8tJExHYWlemTbx2UZ+Xxhz+uTC20GHKDTCE1RMy
22tovror2qok8YKu0LIwfvv9xj1kEg3qImtM90OLGM4MysvZzRkOOskCG5PLZoUq7/+ZtIUmmw5X
3ylCP/aHkc6/MxrX7WBpkxxad6/4gABJ0G0AS4gng29f0LYrKnL22lkm9zblXzJtL7YWSRDCF6pO
Oqsy/8TXu/7mwP75Gta6i68RYeb8VHO0dxrjSUXenCvTab7XSqZOXQ4LM6JNnmaAaXuTK34JV9Y/
du8A1OimnFxWoBJw/PBS9d+uTM5c+OprMnostW3zfc1fDPpwiT6GPQ+cC+CIMFX7GKp8O/6yVu9Q
rrIPm91eeJ/EVarGoyEodMIFm1LEz4ndf0Y3KwZoHfkagdVOSOakm07G3grRKqr042gshHFZyKN+
eOYrB9fv5dYyNPurBYSexnCICN7znQAptAZGmI8sfZx1GU+DFzL6nnJwzikjP/I3F7LrVog4y3vg
M5SUme/TN3rK8ccqyE4e1Jot89OxuLGnJLEARlWQXoBrgmBtDeDx6BIySB/xDm5qyGE9j3gW1yjq
Al0KlZU/wwAv5Q79I1ehEK8ed+qcc3WtKFWK734O+ByoSD10EET4vTSzPDLCiUfxLiZ4IlyssZrK
QD/qUy2b09JFvgeScQ3w3srzIJi37UEiCI+I7T23CtyxHfY4Yt2n5qtFsrrXiqjShwh+Ha3O0Jk+
AVx/DaRNoYCThJFFTBdPOids7tRzh1P88VLXBKcGE4IO8raNjkOlB1J0YBEu6EDItRWhNDUoTvh+
q8/xjAX5RCw4/bQJ0c/6jztBGWzFB5q+sXo+uutY6+tjiYd8qlxMMuBX+Mxvm5Of7cObTz0R+e98
oWIMGgJIyvMMbFtpIb0swu9oQyTy69/0kVdRxM3gx3Wd89hCDF87NuS+2i537CaOmjb3JKRXOTCg
zuVvSpM5qxmnvWkvwUYz+brCIg9IPDEluDXQz8Cj+RSfONHyd5fS+mjpsYiKXqzdBi2mWCmPeA0u
LqlikCqQnHVEHHQbSwVMGVG1pAKdrCk4LvupDQMJjalu1NO5BRxDwQjJKpfF6jcEje49o3bFdjJU
P00lRPPUTd/8HFZJfxHRU504EoEQGae2kmKnxO3A972eMojSODiICQd5UeiNCMdk9adMH20Z/IoP
yavJqBVfb2M8whBcwV92PM+/zf8q36D88sua0Yq3oAMoXmPCA+vWza0bmGRAseyw0z5eKjKfdyeY
9JqPHDkChsjfxhZM/BtjDSCmV4CxsYAfiE51oNtsCT6WzxNwmF2NUTR5W/eCd0NHkwqkx+2ac5xP
HF66DNDN4tyX1ogQjbekvCJsNjnYaUyoVfn9BORwpAlXVLdtea6yA7+1DU3KTtMyKpql+NFYX34m
O1/tji9dl2azggvdLLbHxpiaO7c/YwnekP2hEFsWtrDoqvAB/7iVQ9s0qdDom3YOmz/mMfJDUKXL
9s1epSQQtbvm7qaS2lxwNcmHuKz2vifuTPHPjXvAAtsqER39YRFG0kaeKG2S8g1/Gl2C7STZX4fh
ceLASwy5PcYnGJB71FjjGbM4dCIeKzxTM48Pwqka0cosDcDQoPnWb3tSp8eQFH5d1WoDeInJuhbB
SQHDklvYTZ6TB/eCNN0wk062XL1Q0aw4121fCQDXWQGmZG2ooLQOEFt/9BQWsLuc3yR+YxleCDTF
8kNe/Qi7qkLhyhPzkeKGtl8xCVDICOUuEvFYm93y0XYBau6dvHybopIkiKkDDtVEwg6LIz48NP/S
A4p8Zwne1hL7jYjRLII8l9rmFy+vgP8g75yvwTaQxr5z6UfiHF4Hvgb3cA06McL8ftOpiDSNRef5
UnQp0cudHD6o3uCjpkP80z7JvMEYa9L6fFNliKpfky5wrmCk31+dSI3o4H5G4L1dHBlLaBRopMMo
TlZ7hRva6hNshCr7U/DZhuS0Z6i0OUkOqejsr8ZUP5Va03eb+vCPSbtZcUYdrra+cuUE8xQ3Ft2O
N8CMMDD56/cmJBQvhfRwCHnEqSScCrRbdybmqVejAFXljWcKNZAQPumGlKqnRBsaZji1Gju8dhlO
niqo9bvn+AKfRpDvqvBliHkI0bHc9a3v6e6QuzSfvKOXd+kd3VozPajrqJkHrtfogtsbCdZXEdhU
Dy2kQZfza5KADXU9c0QXThxNJMANvIIIyAB6E+1aHmby5AYD41pDRzT6ZWFC5irT0bpnLQ0KM/ko
9UDXFNl1Iv8TcpqTnrVRu2FV1FPUbpYp0v58FcEANMVXuGuzwlRfju+lJb8dOOp/obk7RRP6u5UW
uIOAVT3YKrwq3j9WKSNL6JmXXwC1JupCJe/EKPxUg9pwxbYULb+jMLaCa0EzcicWRabZWrzBYa5M
Z21Ir/0jQYR+B9Kb06ovcEdEEC+63vXgG/lQCnHmChCPigye68ptEOtF1i/h1VUwoIP00jo1AoKQ
k7vb3eWA3YbyEliuX1YAW5vkPpC2n5SSUH/L+4E3ZHFGyYdvBMZzbqlBFG/ItjdACr0UAnUBgN22
nGRLxRZQWp6LK8cYRQPxB0ksnvRyVTnVTYCmKUHFUMLzni/bFi89J9wxykBBJx1qIMAmOUYt3/uM
Csf+XxGJ4Slm1dPqD/NHT8MZW5EBUJnmnOmW0mUim9fg+i6lSgnZRPB/I+ZSSX3Bi2RnZLsZL92a
NYP8Std4gyapqzoMWQp2XEJb6OGp1Jh3kO1qIFdQ6XVQmMST6L6VSYgbfFjwN2Pso7MxqB6TCVpI
4rY5AmCFV5DQBRNbn6pwLv/+x2wLHPEk5yzw0nIkUVr/7B52/iDRnj1z5iBcezPw7KD/GA8gKy1N
OszaNyliv4PfwvSL00RjbUkrmCQ8nvqFR7EXj7RLqyUZSEdvavYlKLct4P+FfqYBm7geS4RTad7C
0k3zoufnv9MvzALXkK8rQMkPfxOZbMJcxpJeJU0W1UBuF2tEliyEME+0RBOpnx+id2dQ4DUluThb
7uc+iVmQsmuYoLNGwrOiS98pREXo0MsDAnOzqZwVqMzVUjRs5eUQaBXgxLmPiK1j93cENVRpMem2
zsS7Fg0sqayYUTPZkmKMvBH6TW5Ya4v7G8UyVMlPuvmCoHNrn2jYegjOXPP2ehRDafkEKGWo4HWW
/0DFDW8PTe0BfFIQFTLbk1Au7x2SJRluztUtxTWHCCE42D38px/lVhs9Z0tcAoCKF2RBvWQ2Z0Uv
I9Rr8MOPfxxc30ENzNi9+WtARvQ+CUVWrNlQ7Eu6y3hXUMZJ7nJ/mge7LvW2lNG+yLWFHoLtcyMc
U+8u6WuAM2eM3N3mWW8Tbfz4LWoh6jeGh2gk2m3ssXoQ8bgyovi+Ts0P6IOfehbc3RvgXbm8DjnW
zYpKvfV5Zq008D7p/x5p4u4YFuOcVqCN9lb3FMyb1YNXvhN1es6EIyB7rFrf+Onbdm7/95CZ2swP
Iu7owvQfmsO21keBTw9ziPiydUCzmbuIwHv38qPe9MD2C6yfQ2OKAOwolUj5okom6a+wrylqBWtt
Z3873SQmDPiz8ObPUFiN1wTHWkMhrZcBFfZdMaGB8tuKOQqd0ICm8U89nvyKQBkykpmzNAstt2us
Ud94qeb6nc2EG5Zj+EIcEbMld33DhLNpfkJ0QiWt0uGbYwv25MvGlKdP0gRagJWo7W20O2af3nSE
awu9sC5BlorL0udT9PiQJBtliOMtP1Jx1uQb8iFK5EAA7EZKsxX3SyZB36dqFiT3UYU/bKyvFN8U
cjXS7Yxy4dV2m34og0M6soV4iyWEj3tnRONqFuJKbODo531FVp1EzMjJEInyH2XWR/48OiPiwdOF
WwIGXacRcRteBXC7gfukG3ZibpdViuHuLknOV/KWN9gIPAY0hYqe6T+Y0+Np2TZ2sFaOX9B+MuoD
EMZ/q5TT+5KgiL+GG4JinC+DlPjxL9qONi+hAymdEcq4kWDs+CzgbRCzlC/KKDvlpRZD1UwOgdOQ
yIVmYmbGAGuZV3JFUYOIfv/XdLgNnf+h50bPEbCGGFT/HXWhKSEauA45rr8uUtcBGWrhWPwkwqUx
xxFVw65XPVNv4L1qJnrkFXdwutpYz8sD4FWklv+hID/VA6zjbXcSeYORYjcabDv+IxRl8TNrRV88
M7vONkDyJtzSfalh5qHCgfL4UNrWWQlFBNCIiKx7QDi2g8kzWl3jdbt7swDezr7NNAV1L6z/UFaq
c30GVmLx27fRSo4vFeQmTRGO3Kb1ni2KXyl7R6UyyHl2P0C85lvhy93GfPDTzWl123ocJm8u04ri
AGRPkNNnT9RSSSk75ceJt1a0BLIFydZ09xlVwJfaX1X12tUP1DDV7OnklFStQQofN1T8zVs9lvHv
nlDsXRx1EvalAnsurnFDYbUdMw50R4N7aydxZnd+lWy09mrYrFKtOKQEJTLkDX1Hd3EMWMdogmUC
pi5TFGMX2VV0LiSEftLCa386GD+HcGAnoWm1JbL7dXiRKDwxkNZtP9t4S+ZvbOGRrYPJS6eUsq26
WpgAA55mLZaTOze14t7NIq9z/m9OGKC8N2nRMR1/l06pdpRRbsYCgsiatI6uDzqQXnmc7N8d/LZM
tjvrQLGpZSniXyOn5PAyk/BlhEim+yWYdrLI6JhTJxTJqafREEXml2exFp5d9/mhtfCs7sI4e1wS
dFurJ4Oe7pZ4GCMrXL+oCjXtFPRnNaSls4fW/zl5/5c9+DnDVkmQfC0Rb1pPdQf/Lu6y2dJQx1qp
9VKGYeFwlGZ47FCynrKHhkchmQk1YI2UJ1HUbNP9VxXToBMyFM8lgBlDgpiSGxoy0aCUDM78KZDP
UcT2LVkTLrUuVa5375Q2kqN5XeP5R32Hg6ufmQ+kRjOwix8cLmtwzNEGI83qRDzxv7taaaY/LpA4
LqBtlIGOAErsEu3PI35DomPXm3ThKeqQA5xgRKTAo1m4oz0PZLpTeOoNHhZK1yJkNfNYX5x37zaS
fa3uRw6FptyXn1g9WMX8cYT5vGw4C9z/MDpJzIIz0D4T6nG8QiN5Teq3FNR8Imzswud6ZGgGZykz
CoUNiixsJwPZoMlA6vjwX6QQB9GCTdMGY/VPNn4E0OTfe0l1iEyFA/Pyu6YHOIqZSjJ2AjrLKZ5G
ZbhMnTmUxLDro0Qet6YpK9ytGWqOWKeRYl8AMEDDi/xYoyvKe4sLegm/SuDBQUCiaLj1X9IFXcA7
btQ81H9GaKjlsUzqJTJ3o950kCrj69F10o7JPYTJDsCtbYx3niTXav0Ba8i7jVAqKExtgXgZyzTL
MGXlPbssUo/LEd6uJ6ZdBatnYwaGAkSSy9McZSPPyvsypDwdlCoXx3f3x5G0XMnp3G5x52638mg2
kIie//uUJdTgkaXVQi9hPG4pBjLr+hU06ew0BkMVrajMNdNyBoAHnNy7EAfXjGGuQ5u8PnUgKu9v
K5zA0MXnFowwRj3MgrXIHPLxMGQyRSFd7EH0LlO6gu/2K7+fC1R3/DxzedlbamW3iu2ZCa+2JNZu
FvfH/hC/8ItnNbdyClivEbiKBpcoDqoC73V7gfIGNPxGANHFJoALLMgFShd2coMp4oWIp9HpHsmT
x5T85star/A9c7x7G26OCO8fIE/KF4vFJx1zZDkl+ntU7cvhmOk4bAS3VuCVEG/D7Ow4d10Nf2U4
RNbivFypMS1i1w9QLusPfg+nG00DuWcaUydJ1JerJ0SLB6yVRKiK7jAPSLAxvsZxhYVCPqPELfwX
1VqbP4WdXpcNeMQcIjMXnrzbNh1e0Tl3fbZ41U3ouNTqWZkizpxisGLqi0mI59jJITpDA1GafN+x
6hJPOe0FzNtwerR1jeq+5TMPZmT4vvPGoOToxR6+16bHCx2UFgP36D99Zfrbkpolg4HumI7FzMHD
gbRQSjquortH9uyIOc2AC10wUwdjLV3YIsgfpQ8bLgNYZ8gzaRFXdfKvwewcL7HyvGUbwNTQH1wM
SzA/+vuYMmm3QF+c5ELqLhR1lbbVBlG/ikAJt5Ocije22Vung13r6lGxDCMcqZOOfq3vw3u2St4T
NapGYu4LMSdKYqogjv7qCaZOOHnULzNZHfw0QKYrgBGuS7ieeSMCBjzMIsmSqz6YlHWXz4+b0Jpe
yjgBQwrEC5NpZipRHg+2WqDj6UMLLn81FEvWzbD94o4C9WblWlCivkN6IpY/qGHWgrR7n/8EcREP
NWV+JOgJ+PjuBdgRc8M1v/ae52cjzeOW9B4uFV1W5prfkZ6pI0BhCwVAo7wvQM4RTaaWz2kLX83F
+FgKPL5L4PXASQN/aTZma3aYfXvPVGQj43SeiPtg+LEH2/WQr43K/rYX2ppQ8PuXR9r4xdXhUNqz
9SiT6hoAw/mz28UmtrkmaXDW3fsvCporiDi8HSCkdF56Hg8MVKhBaqDtLZ97sjaaOsMZFOOaMZcx
RUdSVGpY1nehcnNcjp3viSOE4uJH3vCu+jYjcHwCLwO8h2fKqwoi/FLrfYrYgr/ljyyvu9/fL+ZS
26nEzUjZAf4DiBU1yhDPKx959tOuZfBjslVP8lS1TnyuE8sCFjxemAreSpzAW8qLbHzuKz+2x8Gy
ulD4DleJjZYbnL8K3pRtC7s8M0L0n7KuHW+LTHR0MMdeEtZrh9/vB0J2fXUkRpKRhhdxGl00tQ9L
S0LCHRv66mfuQYIecL35fW/BC47X8fpO+i4DxLycB0XiuPDpicVeVEzs+UCXvrpxJjE5huoiREqb
QRA7BmEO8cN89Ky2gx87WWy04ZU17wWe18NTASI6Ym2o6+mvNIdyM9xexxHbuLTEIdMk6j8kxk/x
6sRwJNcwNow4Xg/SmNqEdksXCfo7zbf3pcWlFNOMjHlQBQXk/9UpiJ6DNQXJKAhH3RCJ2In3VG/6
2quDf5cUiaANGxOP52cIM/VkXaAc97il9M20Z4GAyzrtftBfwFZf7RJT7iYMyr/16mHCHNyKgYl5
jnK+a/zIqg0PsDXQfhpY/+DZ2DAqwRurlD42lxK3jQIFxnlFFEgRJehalyG7OWdRZSts/P4gKhk9
s88WZdOVf9lKWCP7mKX/5fpYZnP8IawIDmFmqvO//atpijAni2Qy98rhD4XD5UdVNUaO8og0ree6
T2D0oPIHPrQbBwvC2TwN/VA19mDtTNctaDX1bdhGH/hxmL0KwyiIydIicb8dg+TGX2+vW6jUpXU1
GVprcY7h9A5cd2a1PJ4LEsIEKflmtQ4v+O0CQw+slFidtf8ts8EAMDbpKBFATdJh+3CZMnKFrvBp
INxSVjeeZ9rzQqTKH0C6TkPAPKExV52XblH/r6wRLLpkwOgFMWVHmohlzjeK/oZvfomB9eFh1LVF
/GnZGvSJ5T4hWfRgx3LMk1Te/OR7uQTpq/V+YK8Izy4nuws/6qpm2wTIkawZHTLbGuzqHLUAt881
Mcb0BfEJz5/RdKGfmFrm1Pfh8sNHaWC57v5t5ltOzqmWRbuvilu4YxPiHeMlVIEgaYXEFe4iKqd1
ZRkFMOhpkKvBJX3LqujF4YKa8ei1MdE1XFgb+lRQTzADHEp73HlScgSG3SRZOo6Fu+Dh6NMrduAt
+MidyMkd75guUbElnYh73wvU9TUccZJIUNe5DWY7+AOKJD1W1q5Xy/+1cp3vnREfPMuZk8hUrnzM
oNRK0aAIGtcafTE09Fxg2qeRX7ZMfCr8G/nOi8WYRnC8MksVOho5UFiT9NuoTdgkyaX9FNx9sUTn
buD2ERZBKtd6YqG57UVHq6Ql7htQKoWo/fSY0F/ur+MUFwYfOIuPqe9lRG333tMT5Qa7X9QVHVNf
6QHZqKWZIqrYbweoLz1zeq6fdBPU2ufExG2lCl8vOdq5yC8udt99sqo1E2QuaejuDt8yKdAPn23Z
1pkyYHs4CM2ACfWluhEfNCZol51ATq9gPzifRH2LMvu/671cSnh9cIjD8QtnsQQMUOVIohZAdwVs
i1mlbVS1l4MJQZG0p03e05L+7R2IhQnqhjxuqRVDLZz4kp+dSdWvrIm0I2twq8GaJMerc0ANBBmd
p0vEfbzA4RwhWILxG8TArqyms01cP6jhszSymas8yNopyzITnlujjK90TKU5mgSJRhEFKmsiHFjn
bADWJ3/YmT4LsNuRBOY2dbvdC/P+SSbbh94c/VyRB7T6lF38tcDdjYuLDYHh6y2cQa0hrRDxSF3y
5H3FKc3lzIugdRDlp7DsSX76TYtUMjfOtAZ7GxF11K0B5Oz8Td/eHHh2h5HYHg5f7fc6pfNac65M
JjpOD6aeHqlFGkoiFe33iWnzVetOwP2oILiSEK2WI16fDaauRAQV1SYMEC+e3SALw2yPQ3Ejspov
2m6oydR7UdJwLsKZnkF/hGOMGTlj55BVfz6eptoRxVHDYtpNLuOK3DYZFwnRV4tnAXj/UCVYrV60
r+uuVUEnmtOMrmEANfwoa0QSIGctNiWFvRIWllXjVtxRzumvpsMW0ITtU1aqRRAzqFKQyUpcUiwg
ijkGc3UfNsaUMCUag/GcQWrK+o2ZKlOcl1m32dl/Xvs+Nwp8hu/qsnCPizhJD8A925nenO2kPuTE
7Kg+yJyY51bMsPy8O7ngNBv7qudv6F3i5p161mPa/XeQjLcvDgP0nsxnnnw1WpCUr/+uH6/JVxV5
rFvaY1d/yFWRfiakp4+ERshVVOd07CwLNnKDenvEezjui9Zmn+hed3ueESKbJwmoZ/ORGQ2pP155
b5LhNUhNaSGAHyasAncXeR3SEOfFB89QPp/TIdpcOUWTEPDSu3XF7efDhhg8GhN23Sexvhh3tpM8
/d9FPJCHts8c7yTCBWkZeS/YV9fLx4EPssYm826OXtxle42SsyLQMDrdSKLXftzO9MM6iEcYoba5
IS77IyqBi8gKyjV06Po2Nwvade4pREs8e4chKXLOliQCjQZjNGk1KPsrREH99XOuqo6SS7fUQWvp
/kPWHketiZnZPM8ioqK7n7N8z1kML239S89TrvbT0s0nlPUrUbjnIygcRgMTuH+lRwOqpGxcNaT7
fFTQBWcgG8CI6H/dISvIHif/fo8tTYOMJ+HjTRtdhitf3tRXSu/P+GMA6lMxjczawqnc/x+aZqyW
49zrh0Vvn2xixr8O/0veRMMsy7PohGl4M8byI5ed7mhYpa6jgtS+YDKCyy0innj9e6pZObDQAvAH
WAlpVE/MS2tlMbQv9dRfRVgigsaQ+/r8m52nEbZ9mU85LmskMuK7aODH8ZdZdMntYQFRP4I6jdX2
KHqFLHOmeQKYfVSmDpaYhs4oMHZAsW1Lef8zXymCw5Y0w/AGUiJlhgNnAwPUTNy0G8EHXovPzytz
s1C5PTj1xMmld4fGqZPJlVPFpuFcvA8g0i8SLA+Gp/R97yKdsZhCmAk0XCxh5lumaSqG/ozs/5TM
dxSKtdEhbcq8U6xQgTpyeq1d/IgGawkowEJPHa6bC49btEa69vwF88x6AiXs+IagjEImj3QvnnKn
AzXQ5IcC2Wd8Sndne25+j3WBNHIMKQ0026JEYkDxZfA1Q1LZnKNSywV+N1PKPnRu1dJEf/rBpf2u
PK7xaaaPdQ5dSsD+xSLu17uanMVcqQS6zglYkGc72t2cO+QnKl/hEk1rSfvkWlwkkyFDxYKvU2W6
OEM+De8zgrZ0kVc441Jy74c2fbLh8VuTSU73OHgsklFdITgde6MvfQZdVwZrdC+7qNRwlmLqJouD
2C6T3RzFRU0Y+D4tnyN4lDqgaLGDAVAi7L9hrPIq3bs620okS66DasQgdSQYzZVZG16q6mIBZS99
nX6oxylGRJ4gmxjQli2Xk/xpiXfqcH14EgEO1+WXKjiEHqZzvMLr3GLrfJZeZhw7vC3FCOqeazqq
kbGRaEe4R+6ISvXR3v2+AoujVwEa+SFDpk0cBEsN4QWrMEIgZiMtN4J2cIFCXVjA7Q9wMLN3A51Y
Hn7CTPojjllau1JnKq6tj1up9uNOmW8UfVPg6MiTrrGv7FAGfDDAWkusM/aB2vb5nOb6zPlOkjOe
HFJdl1c+xc5/QoAdv4i0Rs6+tHcz+e+g1Q0CfwqcwC1qGs9sw4KKqWzvDigoGb++ln75RMS0rw5a
8Nts0plUgVVO2hgXnTmyZTb29rLZ9I2Xje7zxEvXKpEK66xfmpNLH/EKdBCY4sfUUmlY0WJIZI0G
VSbHMsX0VaCvXjFiXJiD11Is8xwT+zvfZeDyVBgfwVb4x2kxJB2iFSt8WmodkgRhexiTEWQ+cpBK
duqliX6NMxZJoiNvuDshM+SBPm2ewBxbYiFh7rlizkhYCUzxXxvN0pNFDshXSf1nIm30k7Sic7Dx
t3FkwGeJPdxVSDCiFlikg7TKryk53msuofDofW14ldZpMkXBmjcgz9shOeqU2kVdWp+g4OB0qD7k
2I//e4BH9wKYvsKDIzvuzundLJq0ratZu5mJMw/vlBCq/Zwwkwp321ZASJjhKWuWLymXI48hxEC1
vPHoo724WYW09z4Yj1WpAn2oNxFQrTWmZ+KrCx0i4dmwNDSNF5ltipuLBeA2658xXTJ9vbc6ODn7
3lQZHZTCmY9ylQ8g2QSBpZB/EdP2ugefBMCWZ/mjTdSDi05K89U22MlWz3HiEKp78EpJAPKV1HT2
mlGrnjhxDthlfW51cNiVP6rF0cWtNuVUanQ0ZZuSAEtvZ6GYbRYCCGOdl8/RGU83YwtVR5GRN68q
udCIWVIqICSkkd1ZBxfPQXYFiMSDNTtEngkHQTAjQckPLFPxZhgSnixqMJxkuPHMwot8GgJ0j8D7
NGOOWhc3aolHjTvrlcIZmO98sDUxFHRBqfaop5XrFa7dv7sdwa24DvKkNvdyozTFhVb2gQOOxglc
NgTpQ/8eDTjS0n1bC0n/JlI9QhVNgpAp9zpFbZ8XOn05qskHNYLww2x/lF+2tqcEyL457KEpZgPi
wyzzrCbxurDaZ67iB9VQH1Bxqf/NQlGwh3VI/YenIW1gMkZI6ujfPiBkyQV9YTl5RqHeseMV4ISr
BzkSroy6o359nLePRhFtkF7S5hGjmKC3WOk8H5vKCBnZoIJAMWZzATLmdxx5Mklebc1GG5Lb81+t
RTrnlWjDi+3fQidZgsrUFmgzJ/PUa9oAXrRvyMmjdXS37BpZD1LOQgJSIN5K0FrVZmtG7rVd2Jyp
fyGTkC6zQnG3kviJ4BqwTgqySe3w+7GMzmjBG7iWJmCb9xUvkPv6DAH2afwcMU6Vx93tY6Vqget9
Dkpk5SfDDjWjxMyswc92TfSoiQ4v3fEZQMK777G6Pr8prQGBFPJ1eWZH4Mvi/5zb5GC3V92/CerS
DYyaJ0835VcZXkTQyTZaYN+e6PqTO5Zf6XIVY8LmmVH9942j4QmhM6vpoB+cr53Jfqyd3gcZp9o5
kXH5G/7K4cJUkBbncCQmOZ2dvsd5pAeJAZYkgws3dKNW/BzHw3MW9IVwTH7SNyuFA5BUKZy/9c4B
pCsG2hzFHWJn3kE9XliLn3iWHzitybGmU9z4AHfGUQpHM9QDTtTukyncsICR6AtJprL/mPeGb5gT
7ER8HxK+25ZA+AnotpS39BagItdQZlveHL7OSP/fLz+ZvL9UontNjFL8zs0JodrpDor99LLXYeu6
+ozZsoWVmMgMOj11ZfpHW/AmOB9VHebn1t9zpyVhWXhGu1gVm0l1E0KPzCOD1DQI5wfXKiT+uyCt
uS5kCBHICxVN4L1EK1/ZQtL3UiTIt5ml2xEHyoWqAWMWGJl+MjG8akMR/Q8THe/3JXyI8WqQtczI
issLigZoZc5P31ZrY7CeBNrnNPTQaJkTfhOFMXr4iDD5IFj4FiteRu5FTKD6sTvAWE/rGyYv5oEX
CfTdKG6hAtLknWdd8L7ZBlYRVCbOkI75vpPm3SeoJh5emlCZOoZxg2eMumRY56xHPvywjyiOT8pJ
+tKTTJPjCoGyWEQhKtrXHDRc1I9mbgi8lGCyWY5omOZaIFeqQzJzMV7CIL+tsEFxgOPD5DgqxJRh
P2BBTJrHPVPl0R/bCuCqhSUwdAACzBgIGusLfXq6+rmbM4FkQnAv/Mvi2UthwCBOD4PDmec64dwd
KcD3o7Rc1ciGacyLxzDQF1NsTFU9J2lFWa+TN6zMe4IqBpJRnSL4B72XowUdGVVFWFQV8OefpT6j
YGXfbj8z44LEwkKIyqvLGK2ad9bXrE78kha/rZ8S1c10/3fsVCFdKEkppaj3hBzrOOIkJI6nTjnq
jSYLT/bvoUp+UKU2tzHpOQuZilUvA4v51PPqKIZsEv4VF0MwhfRXpjbFPo5VQlCK7lpnddrXK7mf
BJMErLOvUyeWtLtW2Kd8pEI6CARg+7CfglviKDbkfNWitxactuaIyYosKyFahpisUyfyk590dbmz
YrxdTkPUrUHtJAp7YIXOBy5w6JNQu0OqU9JpVusHKooEpPKm4F/b2uS3HH565CmL5WcDeDVh/i6u
fOQcCAFq1WWRczHi7b2ijPX2SLvesZyx2A+u0BDVlDM/lyK0RbxZOgfiyNyNeeLpJhCPSfCuG2d2
l/2HwtODRRzHYmGdnqOGluqLe/a1Jnwm7Rt2WyIf9d3ZtFkApDTcTorYHJDExD+t+YFq9nMeeHcC
TwpMM0GIxIqDOz/wOnr8RuMmIwzUNW7vUmxrps4XzVkrh/rNnmPzV71KHlbR4GSymp5ZjMhgGe6V
jUb5n3Dzr8gSDmbcFeTut9lJdDqLbllMOg3GZx5vXs4SI7JHglVeS7sszQ3GecyQ/14HKj3p6z3Q
K/4428r9akdfaM6+sCmiXZjH4s2Ly/34DACg7HJZvxSLjcU2f6DAETUtNTS2fDgtgWnFMyTtkc6N
rMVkIHUhgSwzANABWoVixdONw70piuLEj2wjk5iL3Cx50b/7iLzHJ0Zen989b2qy4swzRaibFDRh
rnNgPlsTSZYYE9c3abCB9yxTD6zCrkHw45ZdQeznKCnWDoXlfNNL0o/e1AMmth/5qjvxKaFvGI+G
6NR9HvnaEuClL5GG0KjYrCLKJshdo58c3X9VrV4b5wwZC66piNh9KpNGV3DgO4Ma4F87uDhEARq1
Kwnqje4TdPaQ5nFcEwqGV/GxQPyvWJXLe/4v5/2fGk+T6nU/1yB3fsCM5qDPthgM6r2Y9MK/Q5G4
xTOqBDiW1dakiTVQv3SqIbyvOchmAqP+c+QSATa+dLRWuA8QTAZ2GU6qSrd9/aPK1scHS5bhgj1d
a6AIs+QPoaGazQphrLzN1T9FlHua6vpS5Eu8tK55fHS3ywcVINdw759xTF4AqL0bxdoNZMrHqtDJ
sJRQo+mYXXUYthbwxRDgIv4Atz6RiCe5y46AUBFXK0BCV6R5K2SKXNOW0xxLlb0QuQ5iZdFQWVOV
ZJ2ZfzIcUnfWJeb+nVXxr3g6OqHQTOMSdkF4mupVeZPzFvFTEsu3yLi+Y1iYjyybBw9Z4wXQpMxR
uBR/y4gtPjV07/Mb89tnGzDUaQ3DQZ6tO8Ng/GI42FWApG/zMRg/gOQ8X+IyhD6dq6ZjVVJOZc4i
IEqr53Tbokbt6xBit7xLH8xfieCe41tsw6G24kgElyFpF8soxv6YHvKRBgCRdg4MKWRa1MQs8sDg
kdDH2C9JLH77yOF+4w/dTwiusl8J+ook+HJGdQFVf1oC2Prw1S+Z+Fka8blpVeevif8ROlfu7gFn
sZYjqfJGRoR0/4Bomc6dKptjNwfHjL1JunH3SVVL0iJyAiFxajgLYpgQrSU6WV3yoSPCATgnOmRa
7lbUdvavgdpCW39ZC+ORC3I3BoBdch61lYifjLNXfqig0TDHhBnDSpsHHbpIWX/GV+/hmRJFGIZ2
VNPsnN1MwLxmVceqD8qNeEF8Pqki0eqT+biXiM2YxOBd3aYpu7ImvdN1GNLnIWBhdu9X4lm/VJkQ
aO3AHaE5bO/XB0rBacuAWA1/oxNmAT5VLdBhJ2QRlhzEPj3x+zw0HlxHsZ0PFQtNbIuCKJF5RmsG
QJDXp4KfrUWTUTWh0rHJNg8T+RiA3MqBSyNS7tClSf6JdK8omnYt8W3JbBMDnW1vnbs14wUxs1cP
bdIb9Hh9SQ0cDq/gIlCnj3VyXB0YSyCqj6Rs98l66ScOHyddbWN90MxfO5GRxkxUnBm6ntNf0/3W
KRUsxgFFzNVmTnTPSqDXMxd6af2C6lVj/tl1Gqo2ENOD+dW5qsC3RN3E0dMu5G0VWGKBZiAp5r1p
7hJgfmsbkxO6UbFdFzoPuxSvdy9bDm1zIlX3Ici+AcP1RFJRduH0xShPv6FImp3WyKcSC6sS4ME=
`protect end_protected
