`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oBhV/YVloi3p8qQJ0Yy5xcXRamv+6dV8+G8tYeHfUUBVl+coPuMaSBYW2cQVlAxp+IKCvwePrjDt
bSpm2Ptc3g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pf8N0PdJ5QsLhg83hOx4JbFwJyYXijMvvXMDufX22FCbFdaC95vCGarGKA19+ZNtGRXJrtNdqlK7
kmd4mhyF/dlG/8gHRTC/02lKh0TE5yglx7Aa1hbFte0IziW4jYtBQ4DvWubL1XJ+XyqJh1D1/TJH
wwr9V0Ln7Tq46vGbGFE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ehw6fKruSMbZiyplSMl7AAZyELGApImqeXh3lXNDyqfkI4zBIcnEyqUHFZOh6VGK8Clf+w8jEurl
vIZ8P7mAPlvaQSmSl9Ac7Tff2gVUKWDRjL3FWehhf2UwC9zZFcpUUcB9qiTv+6VlabioKJvrYO6v
H9TFiYjaG3y7nt3nbLFks1JCF5kghG89pkseGXDGdw+ns23fc6y5CJG7aeE8pjAj2ZeWMb4c+/rJ
1OLg7b4Qwg3z9FkoikDDK1Hk8MfKMSageZoiBhLKGPgjqw6rkowtH7PrWurRcI/OJ4QbBjcsSQpI
37yWaCsdGOWVjnJu7PJsX1WvSHrFsOdu8bvL1A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oQI91y2ourTVZ25OJHYXW7KU3TmKh1RYWZCi9hrA0cCtEdbhcH9cPjchoa34cGvkYobwXNjOZsP2
DrXuMybb7RGrX7I4W59qoE9cFH968VAPFHG45dEXeXMANP/vxSEKs2XLA+x59B2Bjnbe3B+2oM01
sX25iv08vIJ7EAUz14k=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h/DSZLb0jssOZ/f7BuhvCf97mTFtf0pgXMMrS3xx9yv7a2mkNoxNDytP5EBoGHFHD/2VDQqi9VOC
g4Xa9no+zBE/9vecShG1CWFr6phYloaseZrOmtQAjnCp1vGl1exlrlVBUzxqZnOIOMt8nfBFydxS
wZMyr60i0aErE/iDdFoEFHhqLXUzBVFSEETlobua17+3IFDxm9V4nu9teq7boWtQt/fB3+zIE5c5
gKAur5uNFvY+cy3T6E0+KSw1X+0ixDZuf9lZbo3mAXy5p8sVOejffD48lBQLHLLoRr2TXcKtMwuV
6QTk/TxyDz0gGx69qC0TgUqVQttvYN29R9Duzg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24496)
`protect data_block
4PdNsyTRG0+KCTd8puCxBD+0WqwN5r3qK1gBf3yp4Kj9C/QhK4s1hVMHsc5SPOhqWE4We0mkcTm3
LnDYrzCYfkWyGqnq+PviT74ZwtW9sTqRsomdV4krUz20IIG+xZ8UtX82duTLucmSxipjuE6TO94s
R/7yBqHp1StEtELz1z/3zZa3rkGSR98vDw1e0X8ES21RKFShYMKUtyDXdJZdbE+uw9L/+poPvMd5
K4LBXijhkYfjuBn6Kb3WUUiS3B/okqXIXe1ydveVqLM4gu7R5DFff1gfI7hYOu3eUFzHuMttouLW
9Fzb02xLKus58FwzaFSrafqahoiRDrFRdwt838qLcL0BXgJEQzJzOv9WFcDdaybmYrMJMJvUQVm1
9gHDDLgbWga28vO4IWM8M8gNmzR9pifPh2DZ1A9L0LyC3uB7YOhVyK5T9vZ0OIbM7AtdIgoavrWz
FZ4G5tcDlcY00xv80IeyUQGfq0BldB09eTdhsgW9nPbAILiP4ihJv5ngHX9dx93KkD4QiZyp/yQD
OiVdzQ9THMTwz5J7EcNB2N8djPcVQow7Wh6wbdbOheI4AepjwEjz8kojYZa77s/B5SXnPX6y+tRY
XmDo9dHlW5Pww3CnBeOMmQfNje8upJYcg4TBYYFC7w8l5UcxGAyv5lr/ZHyo3iLVT7N5Miphv5UW
WvzvcOjiRr8tFWZS8dunBIgSLH0PXpYLIKRU3lVD/gjGc00BlbXyeeDHqxEIDSN8nvA9rA8tdeAQ
f9WleI1xEkFZBfrCdGJ3GGEUscVMA/IbdIjYRKO1YXvRDLP0s2BZ1o3trlsHhlc/NcgJngPYXLNs
2EVbVDtwrP3BfwF65y4A7H/jsC2Vb/sw1GgZ3whtjRee2hMoNJgPhw13d4In9UIBEkD68LE0BoYa
KFdtxNBiS6sd9jWS/2qWAEbrhsM4yW7TK4LJYUxbjIHvo8UUUOSbAyKkRzOm0kTTahSAJrcNWSEa
DnXeGMrlVhtnAftnVmkWJBrsr+2uiXwXMgC/xE4tICQWYRB1q5oj2eTQfqGDMneJSDGjuHEZuTu7
A6pbHfPA0r4eGqS1d8lAQZkA/cViN4Ke27S2bQCuKSztNLaezXMKt49q1Kmp0j88ttY2lGWYG0BF
KRoITTtF9BgLIQwmVASloufTQheF9Hk0ZN7+pS9xg86Hcxol4A4doE7X2KDOZ2tDdunCRl41MuZg
FelTXA34efWsaSF/VDgf3XDoFOaksNxo2fZK2bvv0Skd+lf9SO75xq355mj3XJ3s3SSeClsOhv/x
ZNQMIrpBioYOGLUcEMVrFkybqrsiyYA6DhGvZYy7Olxy7YJrqkWdXH8G0AT34oJmYEMc3xG7yzCG
+8JtjJxCHD/1IbZSCBlb5YulDmhBmYtPYSFtQTo/NoaNl06ES2nN6UsMC1TvhgJRrAOoOq3anJ0Y
/ToS6SPcm3aQU1uj/VKOmB8Bo+gFPbUcbnyjwnc1GmDtDks7jFX5tfhF4SbcDJNurXNp8YwxzZfe
qjwgwsADwUhUsMOY7DUM3EIYDcxJ+i3Ytanihh36V0+ya2UVZa3HFA+a6i+vjtTCpQriMCmHCyKP
PsTEy5BeKY2EmC6FQRz/7hEVXKgTYL5ubE43BRi03ukVLvH5CFnV/8Z79tAdDbMlUCyWrCxR04MK
DKudITkzoXdKCHX6O+Jy++BzuXkyzg4FdCFAlcrx4XgIPgipIOt1QLe8CxoddER4aR4wJ4aicXqK
7wqnzOIaLWMl0yXCCbcSJ8hLbq+jpIarZA54WsyBhiycF1fxSa8hUjJLxlxc9T2E4ORXUGhvBFsW
OSQNTFxElGnQDugWqm8+kbbJH0d4C1Xjc7U716i+7WQMpcl7FLO6IYrm9VaNW8m0OlMmSJZH9Y/T
IuQZmGtB3eA4khZ5gbUkPWxer05rzuhltfAsj2xqGD8vs3p9RhrdY+X6MhvXx2rcJS/EmQXLOS1x
PONlvgw1mrzaK3uCmQxb8PsmhLvA6lUE7xDZvUB0zHVYgM/zvURyotymT3warSzrs6W4uyDl9azq
/WU+vEpbPiE/xk4CjdEPOdWnYYzzt4W/xJdMojcw358+DosXvFYP1gKjP1TTVmBhYQjGj5xqgUNq
3c86mqsIZByQkqmWgmwJuObnwSi2xzRnj85808RGQYuhM2sp+adbIuQsmpcOZd3psTYHLQI4qq1q
amdxMXibdxq0DvUH7BL9TYIHv0DPopoAqVruDJf1U7tfh/DVQQg35LL0UGczJa0aqpKPH3iYNEsJ
amhHvYbw5SYE+3E1LPSAIfVMvVmjnHzmkc+8Vhpghbqq38dKR44dt/59BNnXYMhkoZsZbMPtZ4E0
zffl/ka6qKBkDFJF106Hwl2c2+Ht0ALYey7XcsLheGnmjfIxOlObK46Y2ZO+H6UCZpalMDXLgac9
mzHpHl99t96H2OZW/mKNx1xQ7y3Yh30E0ypp1v2hzu2bpqyucSUYsvAzp7T/WqQGI01uP/AoqcPb
ZqEzVyTaM5dOW18xU3VZnYVMHf8zZ6PTPDEhsD7YsihQypTsyObVp0eMww6eK55IRk+FfiuLQah3
vYjyaMgIIfR5uERBBsFf02uQhnXqx4cI7i/xq9/HsjMaZvqApMBmChfs/1+rZbkYSreqP+zP50ll
6Hsf+9ZwP6jmzK8ZsKBFnnQjEWOVBNyd0lCJFLnHD0WXN82gHWjd0s2p+9sL0JVxqvnrNwWsbcgL
2vJQmRsUIWR7Lek7on60qQQkAdqk/VhcKuT+zIZM9HHxmBXxeU7Ib4E/0sySV1I6xdEeGnScdJDF
ukhHzZxeSb1MePMZ0JyIiNYB33wqxfxyk6YF3eKoRd9DsKPp7nTvxRyESo19KP+JFSgcxEgVVdOf
QYYiO5j4To/hLGaZc2VSBJVpbLb2dMr+SESLpXncd/z1JGpe/zQDGc1qJrev1WiCjtvRN5mcv+S6
w4UNmusVA93DQ1k9my+5cTAQv97VE5OH0ZX1Q30kh9ZFCh1x5yZW/pRgizYEzrAor+IHGS1th1Wx
8M076WgQq7K+yN13geQh2DEe+wcfQo+asLuMNCuLugpZA1uTNXQWf6USqynsCtFNq5lOdJJ3Jtnz
IToDwm0ATXRFYTDRldn4bCzhtFwR3ORyROT2t1/2FmITOL3Qhse8kwVyVwwxNZIi1imqWroOo/IU
JLJ2EefaTu25SAMdXWz1nW1+zmkqI7xz/xSsjwmVWU6fS0EJCb5Fjn5LoHqB4eiGzOv3N6f6/iQJ
Wyfjhd7L6WcwolEh3GS0ybjKyJB4I5Mj3WmwfniFbfAw35QnAz7aVMqgktGlVzhXe/8pCkl7Div7
uVhnb3ZCZ5IB2i3lUCrTQ5FKhpxZG2mjAoh8iLohFCVxrUdG1qd3htp5R+QSsXNpluHrEdp0SLWY
qMIKLgRo+XZL6bK5TYXDrw2/80ByGMLCAK1YAs6fz1RFsQQLQHyV1zhZxebLx5dauO1zDbtitF5R
HoNICS4nUOshzFU4sMiQAp9Y6RpkSYVxULIdV/71GS5p1fzUtBxKGW7HJsnESC69yfOe12ynhwd1
JBX2s4cIlowzoeEWQVtc/ObCvyko4+SA0IzDhmpHIp3cbOZYX9xFsf+roqT/kr4IZUaEnp61MckW
vWg/NOAQhXVIw0LBgssLnM4y3vVDpQAT40JzCJNgiJ72qyIzNPF7KgrCLzNHGBaW1kEzbMBOB9lx
czoNepPXyE5IBOiYqSDbLQTWTADgollAq7aFdTgM0INeIc/OJ2jR1d541YW5t6psHJWp7v0d2r9q
XLJBCHqD4KSwnZenSEBMgY92bYAcUYXa+LLCCNW5xFlMajbJ94JnQ8bqkkal7moTQPsNn/eO7jWe
EH3L9uOqyBk6p/IIT44TA2nHzquHK+6KLsxmQc7/9liIxeMFUziSWxs9dQgGj+w/o3u1azaQFN4d
nHE16/lAbpZA3GrDXshrLxar69V7X3pRbW47KXo38W2qASjsi6fwZTFORPal436WZlfwO6hvoVZh
j7bGD45+bFMOc1WZZXO1vmsGS765ZzwdoKptkREPf3327Cp+dwS9YbJcmc4JQuchhzHtItIPP7qg
N8Re5IKiY6tiTYycMInxoU9xgEjGIJYbGfqccAZCtOzQe7u9bXuDvM3VJUDJhiVENdpXXwkhqnHJ
UrWGdmrOphgX4RIPv9cXC4P/dnczqbDrwvWx2PJzwfqI+/0VmhyjgiTxA1LHmXUF7HNt6M+rSigx
vLtC6Nze7EBngWVV3L+eRLjyiJLLgxfvynDjvMklJOwKKD2k9XMBBP7JBXBiOreTmn+T0nB0BLfj
RUxWD4ufr9roNudcBC35IKgqx+tlkQN6SVuDJ0Hf9omI01g+pKS/xk5F7VoePTWzlU9BK2deFwrP
ZtIafj6rZ4zaKJicBCe3EJJeB/yVU3cuq/W4bJ6pS+7wDYHY8axrG44EKYQTDevWb70Gy4i1Yk4F
OtS4oUHu1mU2UCspHP/mMH+1IWrQ2fL3p9yu0co04e25K5t+pSI6FQir88aee49uyS6bA5l2OG24
TVGo8jYDjrRBS8gQXJLavaJUc2uRwHn9EFeUe4zDidgn2Ut2SNGFPnwZEti5oiq743ccW//EKiim
nX1UffRT1KQJmqBptsY0ut4LkG67DQ5ATOhSPemAzl6K92oHawZt6PkpJatfZ/it5jH/Qv3jFgiy
i81UYqS2rxIieZDcPFJrMy7dON/JwG2qW+3Mbl0W+WW5+C/5ky6OTi7GsNDkRMsn1XMI9fJ+g0q3
KIy+la5+c0tyJnzxkVCiGPwjcO2Fc3N+0Ud0AuqNZLU6IXHJG0K975MfEM+o60UhH3E4HUe+hOsV
NRIdvBp6Z+cHG7G9jeMIzjMMfFcTqpvnSnks7NgaqQvTARdyzT2SvNjBhcShnWAQpjdSEA3vVLMC
DWeVwlWd/CNkKwTqXVXAlTIrJx+87LBaqcVeiqGj8B7gBd5kjKGr3E/4XL/B/hxMsXOijVG8qQYB
cNE5l0Iox4NQglpDcdgkII+kYL2stbxRn71zb3xWAWyg8H39JlgWXev3xGnIwp35osbd1NdHj0Kj
yU57kZdby1Pbu8vfhRHdqJemjBiavovHD4mFXzyOP7aekwg/Q84sAncYGFlF/+IOPcO7TtA/wNc9
YbJRHdaIB6Wo9dbU9PyhfuYF5smfUumBUddnD/n2JSk3ng0UqsU6eVjj4N94DXDFVFnuBw+ixa1j
5/LIczD9XpejLXA55XRVn8tgm2Nu7phnwQ7RNfK08kep8CqucYLyT2uenrXlaoUD401KdaEFZNYE
0atPrTZR7Y4pHOw1hbMTRwAwcyYLJLvSy3q95n1rv/qF4NGQYRE2BrqsKz9wwBsb4fLsv0R4fbz/
CJAH5SO21hMaX9GojWz7uqOX2S5PYnNNemFaJ4nyj8y9pmmng+p2E875gnC0f/GvkpdzzSyEcgdS
zKhwVF+1366LKGi0Jc/22fsBIaMp4AByBZqyMn7eC6ygpCchDXC4zZkdCc79HJg9O5MswHhr86vm
GI0apB72s61ed6IXiJadEfrH8/qGqJsX8w8XpJZ2e1X6Dy2FiZwXrSoX2RIsin54Uhr8HjwdOnnt
nEBRRvIEXjFwUExR1Vc97fhdn8m7CZOjSPFKWg/WU1EHW3XfYTbHGEFRKxGDRAyXkZEIW3GDwa2G
eaXEQ0a8mcBluENA8XU0eYqtclLlOUu0UZst6paFg58g58w2XoCMXrYjHgrH2d10I02TzMdEKzT6
hJnu/0SKZbiwNmGvIecEBcLqQkDHt7PDUEPAs03jS3ZZcZBulexm28eU0stHDnRN/9V98lTZdaaP
VuuekJBUgy8S0yWkxYh1tbhAgp5x5dSQym3nlzXYbnKgE7yzx/Cndu6hlZSj+NvUPqPV8hQZkV5u
TWd3r9kM4FZAeDy5Xome+Dj3HIAIYdNr55rLKveFfLZ2Zo0SlsewcAnU9BJ9JRBg5udAHQZutvCJ
hCvGPnCYfF9edjorrOFWrIy0phSinAifZIPiXrsJ7B1M/+feaYDzu+BMq7Sp0srYG3L7EnHoQuCN
xlCdIEeqLM70m0GXkJ7xn9EdxqUc35+77MCKU2JlJznh65mLdzy8ZpyWd67oVw2TeIVNcCwM/3Wl
Pd9dc+TPlWRaV0M96ccI0HwVVMyxoPMA+ihi0W6FpQAdaLbJHtmCeZQB2zMXoe0TLHP0AMcOBBu+
Uix6mG7uGULNtRfDpxdh/5RnwI4n0YsPJEqB0kl3N5kQdqQJe+rKYJcWvu81I/R2cOKLFfkVGi+C
cZRqLpa6xYZ9xuAGefEj5AZriX3fhjvWBBbniMVZW71khN0E2bBR9oUhA444oBYdE+BqBGUfVgyX
742p7dEPt00IAe4LX2w9+e6BNxQfg2lKGR4iO/xXGuGgWl3NrF+oMYNy/uTca+v5KZEId3po8JD9
Gk6FBoJhBnpaxMzWEHQi84PtoEYMkIULCR6+GJKH4VlGSnRxs35kf1aoERU06g6XE9LHJakOy0Mo
5V5s6DodV6fWD+aSnEfHB7RAd80Je/mRMshR71DF/CwxNuqwqsWVat0kQktYSmrT/g9a+uY6YAJ+
o4L+Lr/o57CNt9EtMSoZBaVZvjSQhvBlBkEC8gxiWtoM4k32CnEPkTl4/jTp5Tp/fzeXeG7aEa7t
Dyz0fXHn84K71arms1A3MCC8TTnE91pAm4vLxiRwIkG8phKDoJpXyGQtYKSzVy2G+3EKnWJ9j7oY
+OMfqq35EwQdTpAk4A6RyAnZBTKzwu1MVSzDIpVCUNC7UFxktcSLXZuBsUsOT60lke9AC2ZNugtY
pAozH/A2uTDiJKFHvyHXlx/q+65obnJxy+vCmIimvFh+3jHadityb/Ahn1V1vZW+0rMzPDieMUlZ
QF1eiJ0QmehNgyaF6nq4BYzyoyK6J6xh44IEV4NEPK3zfB2160yNvRjNeWoDoWyMYF6Q1GRBhEX4
XZyQoQVL4c8ilNwWmXi5ESkNZcZ+T6Dcwr3znMjSJ9W8jsjGGNQ2XPxU5CsK1sshJyYPgTn3io1Z
8A5g9T/M/jpL+xL79DOtY3/ojkSU81dNiWGxgwmYsUmaj0f7mAXketb3hKtnijM3LO4w6XMpRLIZ
Coa8cEnhhexZJhFNKqvZT8kAxItU9z6lHrDclpOnfzIYYBd/wlqCr23ZIiSJHrPyFa7pT6mJeRew
U0PWBrxGVm94suVvS3icbAmmiIeAJeCtgY9VLXau27lTgUU8PIf0exlWGvJ8DPyRCLj405MY61W5
5FRuNo2gLK4UuvM+rtxTM5e9rudoY7KAiVrN4FGu6xAi/Fw7vKDACLGgDUFNjJEWiIPUhaiEqsj4
4wRWKLoUzIc/jX+pCyUiltcoAdgkC5DtfZAATlnsVx8jh9B0vbJcBgXdZIzkD/pNsSj4IoedkGq1
AruDzfgk2fgDIO44pRC/i9hItIZrE/HxMAQ6YCslONYdiUfYnQ2jHyhIoTebHJ73QlMfCzDOF+G8
bR9PxwM1zdXrAV+wv5HmEmlM/kR0dPJM8HUPPDLnw3jji8uX1xaw/x9sXyByLt8WP3Ct5KxwklB3
ysQe8NkO+6o97ObAa+d0PTqBsXI0hm8yXMYsWOpjVTRhrZNuodjMdwblkyHpoGIn4dFScJeiWhkT
Xogdb1+jYV+byHg7970UCueSBlBOrnFx+eTKqanEw5GOBkxoFUbqtVGDnGG/hw1anQloN5Kr7vNN
O+JC2Vuw4M3NhXV3xFRTJHXJObzTZqCGjMrQfmbff3qV8KCmyQo74TG4gVXGwNVMM0h2bCYXQS2k
t68C08gFhW7MiDV0WQz1clXoVfc8WZhwW9w8WA6jPLGhoZwB//6H46Ppbrt/y+FgPazmTipQwYmJ
fxBVOh0FJ8R0booHeXTSv3CzCbcPgxs//a+gtS0vyRHyOJZeBCrMsKbfngKRzA6+wRkkD2jKJWd6
SdQFeTr5jD5zQGD302zU+xpMJoA0lHnE7jAgD+LGm8CdjNUWVa6Un6qNihd9nW/8G+c0ChNKZaTu
XJnLtwaaL5wIKlWGVFmCUfgqpLHnrYD0xKG6BxMZJL4ZNHbtvODhIERx30AmIDp22qsX4lLu8bd3
/VnAPiPoPtBca0vQCQLcfiMdgHX8C43Zg9jr1iR2LOfGYo8KTLE9iIgsUydHZPtFADZJYbBS2vFI
L7NsaT4rrHzRvUSybdIbF8PxBY/7xjty2ZHR+OE0jlmx6AHyLruTOembzGwc+ShoVfiQ8CW/lvVX
iJJG76XDgnN3Hbedu7l2J4fXVW0M1bJSPOWs5wnFDtstAnNBCRVdmLtpfmCsEKPFIW3zuO1a4F4T
UCQuWCcTtfY6ZYerirf87w5HplhpPg+QcZONmqtRq5lpBMAkrUxDcbnrTcxBXZ6wsKdF0tJmcLMX
TmrpDwAvqqyh0Jw93+SiGoqWvBNeY2kt44sqFhtruQIA9o6/XJMPZO4+9zmTyDeED87zj7P9eFXN
DeMTyop7/Rltdc+RxWsOenEceWvMdKIWVgBXUY9Moid8NGU7tUqIbo5VOtbExjmnM6T1asAyfiso
O9BXWT9oh284w5SzYueexxb/L5qDBqXTXN+AL0GwlWTTixiDqY+vHSjqdUuVsfxXPtLfWd9VtiJ2
HMzbrgVM2dH4q8qN1XG2viRjU4z4NR5XiLQLIrV3OUqfTeNqEc8PkrzbN8zUmxoYqL0HE0DORfEf
z4hxzCo9i4mPW//EaJI8d4NYkBZLC4dtDH5J8zCr3bH2nTyuCUQc0UIX3fUQyqk35de0yp4xsMW9
rZYg4Qxa8cDjv+nSsaMLDOTGa9Abc3XU6uhcK01hTecSrbhC5JqxVPDaxpqlNlkBgEGQfj9LX8Cf
l/06SjnHtVcyB6p61mYijRyTJ41cD8m59Bay9rHO82pB/EKv/j7G25vWfo1gmCdRRUnHRbCkRhvM
D98NlnDiFlj9qLzhkYAHZ/GOwK9VQjYN5NVeiUFVrIpd5912dANysdat4Ks4uZ3G3aXMJLS9yCGF
PAV0w6SYGpoyuT/UT++id4jY4rcfgn9u8TXjsa/53O5Z/rSVL5IPgJua83y/3czI4P5CZ6PsgXjh
1BebdKNtZAFjmtMBcbzK4QLTiWfcpgCsRBjifiCs2+u+Kzc2s1XEpbOCQ1rOT1Vm5RxG1jc31arH
pw05QW2V4ic5iNuvLGuCoCMHov9FZamGrY90FXkXjE+9OAobAUv+pagPGZn5lmQ0GD3uS7GLduvO
5PtwV2zZgSjJ2cdcAdvr7mjunZwRpIwoPAthMWNDbXzv/Xx3u+RjaOMzS6R/xzodleUA8vi4WEzD
baR0RZMh303kXx0v60cLqatj7b/9U/awRD8BnhVv2LDEAHnOJlEUVfmt6eqkzNQ79V8wUtihlhPF
O9+9sbutI7Oybm6fygQezA9nqi+RABV9/1mFMeuOE/jt8gD6ylnjP9MdwtpHHGQt5Ds/N5DTrjNR
j59m9qfGEtZoKtgLG2kYHppQIswWhcBDALETAFudnncLgeNYsR8UN7g8Q8fuCM+JhL20WAmF2sPx
zt7duRXpR4VOD9wRhg6t95dY57TqVO533zvQGrEsafxgYrJJ6Bk4t7VHx8Ergarp2EziASDhGaBp
NMaWY3WqvAhRRENdw+U5akL8PdAbgeWQPkQgCVF39gSXhZx0LSK2MgXgd7gDBjxL51UPSNRkd3/K
l34pJdK29BLBCWB1U4tHgDsMCjaEWFXqdSI4nudGz8pKk4FzyPWaqGl0vxuE5l3x00vluAvz5k6r
aeq/gUmNqVCxOyeSCQ7aFEfZVbMHOKw/00d6XUAuUjg+567879YsoJZCBAsXfuyErain4QyecbN9
TUbMRCu1v5dfiNCeJQicsd92TIDfnkqLs3aii/FcAuZUDpd3MMgO8BbXHQasXLJc4TPv6nEKcltJ
/5Qc4spdEn/r8yVZ7B+4GPe2KfRM6UZJfeyXDN0TmCahURZe/IaQ35UwkuYphpQEunBHbWUQqUhJ
aBV3Izh0jZexn6bQWDDw7DisXslkG8RcyArvKBwkqHcGzxPnprXLOmcleOJM64I16o2WenzM1TBf
U4ie4QiT/WFuC9G1U4ez/+015P8TTsTijWU88wgQf/9y9btgC73QwZukEWAjpo8/UDwX5h2iW6hD
a+sZ7xuxOxtk2z8urYyHJGWymdgnjqdxOOTuzsdcHzhTv1ErErgZmLgm5KR4RVSOiieGV50n7p4x
IrkL6XiFjYj0ohehf+egJp7uD5j2KAalX/dmHNWucbU2P/XiDRtUDWELFfIdqXDw18R39eUaJurb
UKutm3rhoW2hmfhQ7A7mXSQ+81vJmalwnAGofmZg2yUs/5rGneeAelhd68e+mnhMnhmR6Q2ZBSrw
cDPS8kp2VWv+IikCBHtI2WyUbp8OCwhWvgaK6stQowKxk+gpnepgjsb88yska6DOJ89z0VS6/6xP
OvtQeufGfZpoFKALzdoSEJmkHAiDIRcuNuK3lFRokYAZ/YA1Kgmm3llqEblbvFDDsYZL9RmawdwW
XUE1Is22mvgGYVu3kVAm7SoySmUGdkh2Xn2cJ6Ouw8n9WxEwHvDUEi0ShTFbgLS363baeWFVS7b2
/mjPD9qpdk09y3PbtBfdplSsnPC/rYTh33zQ+qGI668z5wAdbyVwWAgIDy3yoUCsLSZHpLy3oh/l
KKmHkhqV+CGWglaOEqQA8fk5voFyx6zqymschzCEUlL4YM1trJGxoS8UdzIbAGq4vMqVw3jKcBUn
ZJtnIb9YXOjj606yLv5wET0T9LoE8K5tLMiTn0payo8qGG4u2c+Hm/8ejmqWC9NN+zcPMCdphNcp
ZbVWgRLML0Wuv67ChuyAZcjGhL1pAoo7JtjI5VRSGkZk7JmO4jDG1tDcUcs4f/HRu9wEI/zOIZZw
yR1VMVlKm/12UmbFrPfQNbQcHMSCyg/gMNCrkahNMvcrHTB75K7GSi/15wUcvbcap77kyhz8eAKK
nKXXNGXvm2Yx/anyAqKYej50ul4WArvgAWe7eQue5Alb98fXDzAjL6DFc20wunY3EO7wbIoMET6c
tvvuapnS2VzkgJ1+OW7kvJXIWcNpGG0VcNpDa7ZclSEuTDzHWF28ukMQrlbZx8HBpLLnEcKjF4/Z
pZqXQUBcnapl1CUoQo3sRkvCOhhS5aJxmdsK+RHt7EGZKiFA6oLcjPVGhlqwaRe5vWx//eUQzy+F
cYo4DF9WISksbTTwc4MfUdVheWptAW2C9coNDHvjUw+UKT2quO9l0rdJjPqQjOcd0JMJGQwdBNvB
MdqAYX/xkRB0Dw0eS3z1q3hWfCJNjK33jaT72f1MJ+JzJFBr8lbFsunU9lotDO3Dple6VFI2xJWY
ss6XT0hqDh1oFISTDrW+lYc1XpvkB8Xr+QiH0PwA/3K5C2gaZT4LYozHEIZ6SoW0PmUDEE3MFjlv
kjRMyuQSSnWUX1I3dsWrkFY8f4ZxqJjYaUTW/UG69FIMteIxGOpFv3E8Kro74PISJ36C/Xo4nCDH
0YAGmWX/dhbsFpd1i0z+iug9RJW48iXIPrxd1tP6ifq/hzcbhxaV6LvZJv5sh3tlyvT8YpZvVnn9
GbRA9zyeBDAnbAvmrSr9qG2BfWSzil5Nhb5Z6KXX33dh2uEogV+Ov02TyGu5PYiOwMSIicGxpOPL
9nLYsXatHjfeQWg3KNXAyKgNz8XHtlJYnLVaBDpHsCeRFzAeYuRdDXHrmuuq2sYZnYrkHyNHLJF7
f++OmqZcg1MpKJTqIEGG5Gqe9YSYP6rTnXIOlRPTzvf2vUOEYhDI8UGil0TtYn2hny14UopRmajl
AuS2naf3b/Vs6YGnWyPzeaGUUVXliW9bOOcqJL20U3qn6dwORkaCzK7Acj+NqoBPDPOPu/vx2auG
70/cHFCroMEq7rtTa8zQIozDBhuVhSKDlAf5YA0iahoDBRpyPVYunQL3Fva7DXoiylwpoij5OHeO
a5IHH69esSYeGnwnWcyQ9cChc+wCwG3iIpgdANvYW5vlu+JKn5/eCcnZVmN+vC3RfGXUYkmWN5js
4KC6V01JnFpCfFJwtyaXyPS9TYmvH+lSCQW2wtneNrj9EbDcJj0KjjKyrtcXy6yDhrAv15PKVToy
Nb4nzzdibuCcSTlcJq5/d/kAcVs/7DRyEkKQdN+k7NFOfF601lqvI47W3WJWK9DjJX8f+BwDm1JR
whBcrtitHWHtWuMrBpbEylQjZvG0Cq5UkeEF710B6ch5hJ++MqF3mm/bg99uGHh4+667ddi+1Qjk
fSVy8Dj/Sp+tBo/4/08WogJkDvQn2L23QihgYdf3NiAREeotS4X70a5U4jFv0R03rUXSWkfG9EUv
aKfNfiIG1QHBTcohrUdzXT0GVVHHW6VKLOGO0y/PIUWgbTYdzPLBuTJeJuAggLjsFPFU6FEwpYtt
+yRACDTqtI0Pze/bKCL93SA9wvn/JUA5m5YG4jBadSA0XtEk2IR32qxkc4ZK9H7CQhhmozYuTF/I
9Qa+NpSFh2kBuKqmuo67bzXYuWGV8UeT3aijyGw327cvry1Gprs5xHOYZEtanwKUrvGNs4+SlEZE
UHQ6WKTzzYonKx9QIa65ICCFNcb4tdTF92fLl4OW7Dqvuxb8JDX4XGn6BkMY+8h8jm9XcCxnq+72
6pdH906xWnHoretxtEs7E0ghk2sggbMgl/daRaEja2oZ7M4zc/Sjhxsy4ceKD/2H7ORk4vgbzIAt
oH2mI0lnusM9tSAqqX6mImD7Ig4VKwIHKFBPFrC6Csj09GpB3OJzrR4/qJR1NeFc9Q1Gx78xjYhk
yfm1P++VfjGuSSubxUuqrqFoqfs0SFb7UKvzc8BuEh8akoB1baH7+nbjwN+VnrfhpmguqSU2DuyW
jbBRywdHqwVRoXGH1Dd+y+rv3/yC2C8tQ+PBZnd291v8fhx0bcTwIh3G63BX8fAzLUTcJ4GRPKDL
BjnMBXUuYSxYRnvdAUEn0nKwa4bALuoQm9cKAWApa0klLyxBf84cI26w8vwvsq5JiXELHZi9iU01
7bBcBsJhXCKuP0trl3e2yhpeEu0DdQ+QSUnG5+qcm5gUbNzpsgo/5BGwdeS4eUrjnHdk+vlea0bb
cmW6KwyEjq0w5UNCB2ojuKljWxSOATwMT8XrbtaEdgrxJSTtwl9epu8CAox3N6E/2ajz/urGp4Mk
MYKKXgcD7DTEHLE/8LhINnqdTtSAo4XCdsdhFB6d5F1EKjHtGL3ejkQmBCbiQEMN2RmFYv29Gs9n
BONIoMXp5vNr2da1+j83RFaLxDk44th7e2BRQdkEMc/yQ3+R737vqoEcV8RRyrEKzcstnLy4f0V9
Ke9e1I03BEEy7pkMYmJQvW7DcdG2uNj5z3aDBNrDCRNPjtcMPw4WXG8Ki9qK1qXxt3AfY2wtwxBg
HksUKxwaQ+SFTRIFx2CSjlVb5s5J2rEOVa1lN9/3xtn/33Qv8bn4A1RNbXXLUMilBfPwl0LHxDL3
ATuo/SYU6YkVIzOOo+pjT5t6rYBJfN8kCrS3+A/BC4OWg73n1xArIMDU2VgmduNTJ5TR8Jg4KmmV
yr+NIboPcvNcZibZ7ccgO0nlGP6e7MCu98pNvBEHIhGxW/M04tKni5bif55aLgxklTrATSmF8oSY
4i8tOVhQR68V+p2aLi/XWZPtOS9lf8ydgbUi+jq+X4WTdDzUtIQL1u/CWj/owaVC7wTAyihJNnhq
boiy/qqcZL34RJ2nNjCko7juCokc1wugu9mj/aFpqQS6q/2dVjn05Yxx5n3xC1GLTaIcQx0LKO4c
A71XD/CYOX5WJ0hqpefXlz+cL5tvqM2l9flu2EGKF7ioS2Z9dLPjmqfZ2ffUgPlgBXrhDSbXW2Rk
PEs+vFH2afNxZ9Tz0g6gW+FyZKkAJh7Me1xtWIgppiieWGaK7MaNtLBKAvGpLm03rcR59QC8Sl19
TpDaJ/4y2Ztd53DbIRiofqsQKuoUGsHsAeKoLGM+G6H7qn+c+ExFoQBf63GBZnnltom/qP0ldWjS
QHKWnPMJgtQO8VzgZaTMnEipMSEdwLlacoaeA5LqH6REoiemlPMdv70/5HLHMKmy6kuwq53f/XGN
qU8q6as+ENRn2rsjdyZFuWxq+RKwIUIvadxROD84tiYsXWYyXggYxhLAJA4C+6WVnmvUBPKxaxc7
GkfbNNmWWJSBbMN0sufVap7dM95sjRWPP9aY6edz6kH0eNOVUqT/0Og0GK0x/52tjFooCuf1D+/u
yZdh4YBW1o8x42HukDJxpKFvzaHkWF6toacXuHlh06baDOc9xlS2ZgDzJL6OFagGwOv+MPqNjPgH
hVtwQjhM+v+K0FHz+AcjgG1XO4AcsTBZ1JhYg+Jo79qmPcifFuk/YUIkMh0NtUP1Eb5WcfPoVwCM
r3fEFsbgSrL45p/WhE1I+40zYKWEUNUlafS8kHRI7+7TGD2dhHEuNKjY8APLUrgGxjA/XY9qNl7H
202d0Iezy/xgjEo6QBc+l1Nb3lC3lGO6gmRYy7UerG0USmOvYac/T590V0U0nwQsWrkS5hffz6Ky
ZN7l4QRwRxwh+d5b7Sbz/65Zj8N1gAC5ZLBKHwCRBuxlt9MYPmw4eF4XB6IRbXpJD+Mlbivg1/ED
Gnlqb2mtEwfhl/eoHV4NDeuqOuKSFKb62/4J2zXZhmWFIsVieNLQQQ0iK0iSZtel09ivhbkbRMIc
invtCCCngpc3z8YFzPvlhq6mMV+fhM+FrO+lQq0ddLV97T/5ZZAIHH0Z3HFxqc+ZajmjirThIGWm
eW/DtWLZsgorJYQ0ghjioC13yvRL+ov5FgyiQOjWPb6DzfJT2VppgVozcvwconq1lWh1ViGawhMB
wREHnSYsjZTbApp+GwySRnroK+O3GubzYhN20G/lr2heLQcshgSmvGt/4CrgQtByUSl5HqPWXQvL
QWCdvp+GcXch4YT9hypQ4pu3qmw0KkmtDC7O0pfakNUYdnI3Y59T4YJwKsaMLH8wZ5LyO4c2mIwE
q65rJ1ewocRXjXbsspNrsXkZQqAyiRTvZk7nBg0awB/DaD6gDKNeImTcHuLDO6Tyg15hbiz6ugHM
1xaKwe6KbC6WiBwu9yYaQqOoXIsOlmAk3tLONKZZHT8yQchvrcCzd2QsoWRTOQ3kdSV1Zycn88w6
EQDcetv62gJVeR/IJga06PnEeH+AWEz+wt1Db56qxZQxrcfQLQaWRRWhYvoj4QNGmhFx/K9JutcB
Klqisx2ns8BVXpZ0mfemT4ypJniWMedTlGE6opzRFakAkuvUrT2ZsL0p7ML3ltvPvryEkrfwbSRE
bSiK7lYpyQ6WF29AcWkvycAi9oyl56ii0Ljn2dzzrMdFdmXNaj/VGiPEbCqIcN/lb1wRI1EPmrXF
x6DRz+MROorauZv9xHRSWR4jthyJyTErMUHykv0A1AfvEVjyyZtHUUbbWzEV5wnrNiyAuZT23OXA
BET9o0egSg7l858gsgGZiXcdwfGiDbpoVQBdFUuCOiLVJGGhuYb9W0VmQzqo9m9lnpon7+9MFrfz
vMXTeSoTdoy3e1i9QKCYOPwuGNAJ4bsXOQlkEMV005/lCDCjXTvutBR/gPfInIYJTH7XYur1E5NJ
NmBYLPzkVgHD5EMEGNt1pE7O0fWSOANB2nS/l+Y5JjMCtQmduSwVKsW0fNaopRD+MRMB7DUU6gKj
BIFKU0Wz/z0nnWGboOWXd3UWcJI0/Lc/qbm10Ao5D0v5ltpsiic7PiyDovHVPo6G9b4FpAlRE5hD
HebM3GWzr78HRAdZO4KeqCtwanWDAbRAZKGe5wRUzw28Vf28sTUZ734L21TDW53knHTTPeVxeK7z
Z506v9cBYncXF44kS6QO7/65rNSFIUmg6tNoZf5y8vTziBWPGXIe9qezdPOmQFvsJ2EAvH74QN01
TnpMyJBOv9itTpeCTuMpW4Ohy0JP904YmbHgnGAlWD4G0aNX7TK+gZe1SHI10sFoOVcWtbE5drPH
KL39JLO5YkWyFORFSP3kRD2ofRXg8wwb7OHle4Ec8C65AYrqEo/8j1Rck+o8Gfefu7uyZZxcEwH7
IVsfHfoeoM1vijPBjLahLL0AQR6H30Q/HgYUfqkzgDaYJuWZ4lgXmM1R0g5peg2n66qTXhZjbgLX
BwhD0Ey7k/1gmVTZua+/ETjGevQJeGYswRwvZ8nFOk6Uu16Nh8lG13R3+eOawtfiQC9WIcY7q3JM
yRu9h/P+tfMjfKgnMuhzKG18HO7PozNaxjnMQqmKWwsDvlLYTxpQWeafbJqmAmvQs1j9thgayL3+
JafLQXIrA3hiQ6viOlVgBZw6RbSTCxv04HHgaEO/zWZtFM6zLeYliXUQysB71kytAKzn5q1NnoWV
wpUROi4caKMAoXqqfqg7poUfx/VtLsN6qadPNgJNTu3X7ZZNqHOQU3cISRT2HcS7QZAdYnykw0QU
yI35loQq4DHcyBbxhEnLGCEntzej2qyVXIah0ERthSkh+I4F2maxWSMKDZuHJYX7JT+zuOv0/7Mb
4HARxDBLLf5Hld6T+Pf/xcvCXqyyF1gBnbd+LMEDWbd9WIMmkj8wSc/+Wf/vMv5xeqpJ2SgGnSO6
L/PhszJMtBjxmdcfzTlTWQfPcrG6aCJlZNpsphD4CQ8SiHNdCTozn5tXQdjEHD+rLryEM/4H48kT
HTH1pSUt7C7C61UVe/NVjdIFpVBEuM9gQ9njH4cSsgWkMmudt3mLLHp7b79as5YiFfOLIpQPnrVr
VYm/ZlMijKUXMyp41rdiwP9soxskW1+NAUXLK09F3N/A/lRfTM9BMKzV3mllO2NKJKVCDrxNrE7Q
ACFA8F3Bsla2WXXfvOpHmlLXs0UiaaiyHd/vxuTFVvNPXfRZeNiRzXJVCk3EySAKadVzldtdifqp
srQ2TsgWImOsRGrFC5vLZ46ze1EJ7bSy9gkeqEViEEMPe2gqB9/CkLhrOXMD2tAw9KmzvARFYgX+
0N/bpE+WHxnEitcPWlphZPweHeiVrMMe0FFxMyRjLe5GtGpxl2t3WUrCUnfuJ/AuTqbVVAobWhd1
yy4dNl6F9gaQKpO5keg3Bp2MHVjsFlH1a56/kEsX5GrtC485k+kWjlNJZZITI7//XViim0sadAyQ
Ekw+RViL6+89/tCCMFwulso8/rYQM/2VstaLcva0KXMrX7TRrTTnP/5jpanFdYybJK6HnvNmEe5g
wxKzo7CD4X1bHzjR20nxxltp1W53jZCWQ11UtbBbVjMHB7rZS73PkWA7o2Y0R2nBaieOXIKdTYzf
Pvsl9On3vVh8nca8FkS0WNLq8ZRBXpmaP2IOj8R77ewA4CH29zfBryO7BFxw4e54G/1jeO/SGNoq
F8oG7YVSgt3cG6+blznIONDYoNIyuCV2P8sg+g1LuIn5QEvY/qw7aouyU2mt31WhOfm3u9tIzZBK
dIDOVvPYM6wbEYf093Q8eDIvYejg79N1pOck4CkntOWKDaIPdBOW829YlMF+kOgjpaBxoUg4RZjz
0GhdNUtfIGZkSzIUcynYhQkvC/m4nCvou3nuFZklk9SMqlqd5GDgEpz/1YUZibGUPhgdrlVpkiai
4K3hZtHgh0PhVoxU1qhjcYfaxT+euolAgC2rgfKnOD4VxcjY+AqnQel3VEadL8suPxzNaW1zM3oD
sXlORXlssnBWtNQzBrloKtSid+Kf1DHVYHIlzAXbdlSJlEpHidH5/QgBYIGqhiNy8jKXGW8VKQ1o
QfcxJG3J1QtkFUaak9qBcxFmyr9tFxR/zcbGXPu5kUd73ygQd/xiYGb9n6IOjmddUBAhxL8kN5EM
V2JpMblmubacGjX6yj7PXcXKMmiG68PPyYstAp67VCmb/Ix7+kxLW341lsCG93lUFtrusxH5kUng
L7bbt44duenhwhhg/TXOI/IHpWjiVW2zMj3FZaWgLGxCdlO2XrACfrceBZ7fiZHjLTAEM8+Sh5vn
+rgCtac/BSw0qTwMwId8nmd1iJ7dWrzMyWPnJEmc8pVmeBN3cxQ2yXa3xTseD4oHPdQYV5WrE4AF
1YHIfFlUuu+OgroSsUyy9zwrZuwpU75yltWQrPuQk9YZiz8LotEJ1iDiDl8xFv3vgoDDw96MBAx4
SWKBZjx6DY/CX13gTqupc4BsE1eQboWYzjcePGoqOtP59Jf/y9tgy9zXnOzFmtAKtA3R7ANXrbXW
6S6sj+xp11J3bv463sHP5LBbLE7zjfZtTkACJSSGVXdeaPeBXEN0iPnEyKcyL9NYMZe8qqlHlMEo
z/jxRMikAPsrbmpH7pmoBBTw/93M1ExVVRIjhczIdasednCSK9dfQ+Byd6qw2CWWzORswUVV+iee
gUooUJPjW1H3j1ySBkEfBRMyBKvbLeL2EYYCHKE7Wh73m83IndtB4nF7hDKivgFp8h4s4dgLIAwz
nqKS2AKLHq1gPPfHQTxb84ehtg6eqmpr50iDbRjb6vfDbvfWKF2QwvsvhlcLKW4JXzTfYKhFcRj2
e4jdjcnyCe1XkID71sJMvb7tb7PpqaY2tpe+OhDhrOJUdsVHEvsFU2ADhqG6d2rr9ZWEnVl9Up7A
86koMUWG2IEk1v2mrLq2RwjmjfaPC5i1vsp3IMRzv+Qvn/UH/pC6euwhAjboE4jhV1TCMrHxC5Aj
w0JRzbCuml2m8X90KOxuYUw0/2Q8zCjD9ITWOe/TfbRVdgLL8EbY826Qb4sTdnvGi4ex7Bsl/2/c
CCsnZeoXYsdm/0tONlbkleA0ez5bpfSEyqsPwYFW9qE6jT8l7MD/l7cMkmwEXLiTkSyx2qx6MIv2
vw4bMPxMgcv8/efI+7ijYN11GPIuMdIoz4m2yQHPK36JAjR7ToUZ9Wu//D9h+qKB0pa4EXV4J7pM
VdYfT4yLrzwzg4tZTYkRxdXCt9BL0yFoNE1y18TvL/xllbY/UUWjUbVxwjblOcbXshtH8tmKNrrl
+FBZJy1YtzGAHbwo6BZTOpbTqyLrZxTFbXtQZ5MZyztuF3UN6gbhFRgW+3fGqzyBUMk1Tjru1Una
o4+YpNfUdqzSV3GA9ng9gLZDRx/r3V4rvHM/MwBJHVwt6GSb+g813Og9Ahr6nQyJeYrxWn86tBVj
Y1geai6iDNMYC+KLjN4SAWAb8EhEpFHjBR5NWp0jl4Dd3psJMxA6bTHINRY/F9U+SF4bQIhkOMRf
6+klJAooyflM35H65IdhLiHg7lrH9pqf8ICPZUMxELp8VM01lqf2H5R8YgPjO9z/y7b6UZoIX1KU
nh4cPNkhdrsUonzxh+5kI/pDFk3iUMFZ5rFK0zlKqDvQrAoUocaD1ewiE9ONfGog8cvFgJuucNdm
epMYQuJJN+D2goEgO0J2HEDDoyOMKfQToiKDRxguOf/HwiV5ldMW5NaBEknWu3U5AMtROAeI/DiB
kVNy7KIfFdNdQTryzaRuLNMV/sUc/9mN/vv184yQla679KgaFVk9YvOFpq+HtUUe/aKzFEWTapCj
n7DHoQYddTPIpX8Gpvof69atbTzqKWRgdicNzaK1m+wByUeIKSG+sbPQsWuofpmo4sNbYowjlgDY
T12gkj47eQ2KxoUawbuvsx25UWA4NfxSDFPZ7qSMhAqFtoOvvkGwoQ69Z0nHcP39ZrX5qVnmDloZ
rCEPXPPDUpRaf53tG+3YsCnvIltt/o+Odlgq8RPf5H4lBlAPYAbqEM6j8GY8+AvRFTsiyZY8dbdf
KbTj4Rx4K3boluZvsbENisV5Cl/C2aeeqiX8LagvXfKrYWhgbum8qEBZjs6zFWnn/EWROlET5hP3
WAqTgRJurPXMnCXf8RTYb1MWky1sAlHY0H3qHuXj+EZcW5jg0fdDCj6AuTbLbzuuqJZKXqlktYb8
yRgMqev/KchMWDYkOwj9IyRm3JJ0Cuq5D4b/TiAz8bISNGBMNscwS8VkOZaUncXKYyPNkgMlVGSB
Vg3lz8Jdwp2wM4S97cfmokV/aG8nB73C9FfaiPyfa1NzoYXReWYt7Ud1qR9hoproWfm1Pcn/cbum
fwYPPFhTf7PMqVuW7kKKADoJxyZ/oluFvVxYCffVx+uH+LSwzvc+Bx+UwZwCbttCIkZY0X1kCPRK
zC1YpxN42ZvweoARZeQAMtxiffYFAUwSGNrAvuV1FVqrX+hZdvABgzc/YsuE9tCPEx9NG3zNLaND
xSTUmlW7Ka3BJJHXMzsWUpxpEoleIl4sHL9CYy1s6mTq9JYD0/8a9ikpBeL6P/k9S9dK0JPS9g8Q
0jwbKk7PanwMV8hpiTQNMwvCEorinA1UvphoewJ2Xt0eHnAwQaWOE+2Z2EBNuePFHlj3bdx33fi7
7QuibAyaQMiBIJvaFZbBLX+tT3qXtJxDQ4OBpbjnleqNs1mLz8J7ylFZyFDcNfp6w5yRMR672qyF
DWtNIckcYnGtJvE5JbeLSv4cIqWvF6Ve460dVeu7CnVsR+LuGIIzfcYF12n3+xwlf3UQq5hyNOaJ
QxaFpCPfOim9J2T4LXVToUb7yYCVVB2kOEull6sbhCgE+RBZkbMpeL+LRfA7YrG83QqNNKnr+aAC
YtYbJzrIcy1LtAqidXoqsHtgWGptilbbIGaMvroEojdS9DlOKmz5reEYOJTd4RGNPsYfEmnPqvY1
DFR/J4DDysEIhIdySQyJe0beS9XQwRSHzGlNQ6uSffH8bpvnSPmqz27T3TA6v6jiHexChNGeJi3V
Hu1g//n2K7R2eZX/+41wErpJIW7zp2Sw667Qt8lYCCDU2WkNBQxElHJUHN8JwpJaxAIa94TiHM1A
YTXpSISsaaJPVP1+KZ0n4N18uyv8zM/1snxDH4AdeKJWrzqx04bBFRjydbiD3DB46pw923ey/zcU
3eUg2aYeA9xW+RrPG799OUNweJyiAEtxQA/SBDgBm2ibqxoeAqAGK3x84vZYJYQVr7dqaa3uraPT
Cbvdlu6xDbxIObeG1p30GeDFe3mjzPYf+gUYjD61TRJZqxyoV4HdC01ovf+8lnzUpD4EkuPw2kwW
+nLU6ambC4J5OajJoC4auFMdqs2Re5a9Q9bYNZxiWhHJRTjerRFXzbGmRYyUfd1xpybd5CkhbLjF
C8HhY7A1IieLflRcp9/xlZwbrUeFpaMNNtDk4/vzwoAGWIhzJ/xLzR8kw+SAagP3mUcD0wrfSVBd
EkrfQaavIrR1Y/sXBMXgYYEIvotT/KqX0zOoJVpElglzk9beRmjfyYHKedvq83VL7xpqwNElv4Fo
zWoeBWVRrYG7JMNYwvl+XCou4VicfUg20ljQ+uZVlZbk1leRPTxj9x22gZvKa4qryOM25MLwi92M
sIOoZUlvxpChQarSIvKzWnS0wWy0ebYmkrupy3YnlCki6haakSvNeHeKWyyYP4HdaxeyhBYmzWnI
eHLUcHQEAqrU9HzSc7Kw35kRlCNn15VBvMaTJEz9M1Ir+wt5lnGcRE4D7uTuzNX+r0rgjXuIYl6h
f4HXtN+k8lbhSUpqeYQH3Tn7UMEGjnOkWWiFHN2xvuvFL6VgHu20X3C7XFyMpBUxG0J0yJqklGru
uF/xnczeUrXSr65VqueRxQxsF7AKzi456SqbMTMu12wwxXUqAtNyuCFv+qJ2MCi4KUW0c4ZgnrIF
hVORlqXpAGQXUvlER/dGvnrtVI+U1ZAAFyZ2MInNCwQBF8U0SkrLiBlpMXueiyw7Hbt8y+gyGAcg
7l+3q9GX7tfep9dEd1GHB/s2jAGC/nd4v6mIrnDU/j4RTIN4Yueqq6crhnnzTeMym/rLv87s+Ucy
m6qh+lKgGfE7deaxIJzaeGiMsc/03WXNBRD8g9e3wTZ/lBMXJhroLHvqa2bU+VJJadw5olt1dRrW
iJ377KXUj37j+uj1bT/r0pmAHJDwsvgov06aRCyspEUf/WaWcO2y4s/BTRP7bS0BhP0tsSsmFLcT
HkcQ7j6YOKgHo/47lG6I5ktzvM1WwZJ+DR+JrVTb+paUf5fGwokt7AxQU4vjHrZgFeMFlBawehEH
6CLG9C78IQAZ7Il20lvxcP998Gn2bFV7gTnMb5zOcNa8pMp8fWGNo1E1lnS4DpsizaEMjpc3TMSW
jzUtCGpST3AHLxBW1dPi286jFk4kHVe1na29kaxwRpyHL5KNrLZvrgg/j2ika/UHdjuo3mqP9aHO
nDoRany0xhCMAjFpldV5iqqWiSUTickMI8wrRLN+HUKGT2mBY2KhEMK7SCiIbQnfZFo9CejjW8vw
picoTRSauJ9gKa67P2Jp+LGsdIMD8lwwYBZcLURW26d7lKgsPVWRaRzrsgIqJFau1Hk55d0ibJ6I
utL5O5InFWDdGHo2rYEa/xgDpIjqcySMZEiZ0yTaic/ms7hMayskxin0NpBq216YFqARoNIXWWUq
INFQEwmt1GNcmU8sl8dic3cQG0e43D7c0W8MYUkV3jK7gwFhupnBaSBIEI1I4ppQbQx5ZF2QTaOP
fcdo9KEkc0BraFrurXtROpl+UM6YX3bZ1HQQ+2rS89/7bicfR2ABlwhImSIantJIdpVWZ59pT6wL
IJ5rOnnIudLP4ZwxA+TDTmMqDyB7Di+1zI0JpE+dXvkHvBx5ExVUXzHXkchi2pulFP6FFhrGfK9d
sGyxpBat6SLFu6LRHglGXrhyMXBl4nD9pbfZCxAEHcjysyKFWEiGcoPZOstVbsla6Fqm9lm16nLL
BsM5brojanbMkfb/v6G3o9AsifynKDxdFuQ3UfXlWDBzSLSV6fsdCTg6lPJPGz2YSJcHx8a5tdox
p6ttZjMWZBS0e+4SV1WnnFiIKgs3mlaREXkf+RqRdvkAjXP2GxfiHYuFIIqlTjnlgik9tKpIv90r
8D1b9GrIJtlTMl7ZhcH6dc0egIluY0TsZo/Axzd4w4er7Khgbif/4gP3C5/n5LYKKQPCUk9e6Pws
CaHlQfcsOAiFpc5+cQeQ0zWJqzJy6xBYBM9ZIscJWCzulBRoSgSf6czvJXsHewR1QxVBJGtVn2/u
l7AF05RHxYrv8D+pDj3zeyEvkP+3z0lxEZNodu+WV7YQpllEOKtiKiCzpktoP/PxHac52VEAt1xC
j9Ur6jPcYW0OyG6ovwDWdSDj0wYGRLPIIPRE0HRHjOpeQTmJ4xoUtUpn5L8h5wXoXHyo3pJP4Wyi
L4WIgQHzDA64pgSBfUP31F7xEO2Tx7BEu7wAiWoz/uK2aRO8zKOu5wIUNWwdG4Rd2wBcmMIDdOEa
ekfI6HtuWUHpVwr7lyTx+Z9oMw+8Cooa+57IdG5McySfoxXP3CHq6kSZaKdNY9VtnH3g+FeQb9t7
QZDpFwGe4hNH0VPga3/o4GhwwrJgliaw5SjmZmwJ9eb3WrFNzBVF6CFd9brYRF+FK201AIWalDY+
DI3btaWkgRMLh4XlrwycFZiBiRFpBrp9I7TOjFBTbJAMpbZkiEHmat8nMSoOlETx0TEslDTceG//
WB13tcfqWDKu7yEAV82ZRi9vNnkp6NdiS3TUnPlJpvTm3oPXD1k/qMgBkLhj2wcKKuMtZCUdlWIp
gw/eo8gTYyKLI56YZm1L5SUM/0aYjFIym0kjAaxYrEbO/8zGxvSgH1O5fil19nGjvH3I1laRqZKx
So3ExK4XHcI6I8S3c8QrgO1ZyOX7HeZLrCHBcjP2a5PIzhls1ewyS/gkSdiajrIPhilgYs4zIqJH
61r2/VOHLz6oJl6Ysu0elNJhsADGG/045oGzIOHgo9n7KO872TE0gI8CgtKOM5jzCTcoUVp9L+Df
f20/qf9fKUA8ZWK4F9HLUWRO7n3fkrxsT0uhf1RCWA3ln2P2i5hbeyTw+eApuiI+aNMW0xoZFHnx
0DO9n30wvKoXPe7MdSmiBogH+waOEHUvhjFxlmy3GUoKl5fVV2rSI8oOvoYEPHkGnCfwE1oOPjA0
Z4DJ3vI9jhpIaMYrdI6RtquCUdRBZKlWr28JyNQQeCqmCW/lquvLndv4K4eVEdEIwuRM0mVO03MV
BB1JFKyTPBmpevp4DKPr3mV7nXNRCri/PWch39XM7cBLFo9ngtaHHj/Alef0zLxUioNN5pTmbRcu
ElzaMij0po7gItb1zMTgmmvHgTrkpDxryudWU9PAVInDd+DVSypyGFhltozs2lBl0gVqv2OM3JGz
Z9KkIKEU/0jrrth3n8Lq+PQ48ugCkP/zK0zQ4uES+XxuX+7tiflMHBATADA+aAGkwDR42w+dOtPS
yNbfmQwZKo3lwvP6VwzB9IW+e+XubQhJG48nhtogwztVXcvlVrwshw2S8OUR6iIaV81AXvkM+CiU
OCn73cdKgeP+92uvU6oRwBCd4SMqLL5bcqWeYkvuyt5KD5EzIPxKTqW23qcrwTt45rOBqDTzuqlD
MSR73IOTVp/9A5OMGHtv7ctJUh8HcDqSvcQ33uiJ1m0MIj+Y63HmCyxO7Gm2W6Dg8Gf3HQ7A0USH
nvEO6W5Dh0whIlKGPyTngW7nZn37l0S1b1rfeH80LpUQ9/vlm877HGx9JCGzc2tX4FrYSmohSpzA
zzy6EbzpzUQbs91Ga7f3+zVRgM8DnvAUkdz5/gpJ8b9jzRtFBIdrvg0cGTEXi8HUokHDGqys746A
Kpo862N+YxLlISbLT6dIPftSEue9mqmAKP3Za8OH4dw6FHA1iEMqpMLbJGnT2ZBm7fsUpinF0tWc
/xEAWwy0050OmMzbNMaYgMIYEk0v+YajSk7HGr5DICf3U5yKHoOm+/mql/1sbr6ZTj4lyeX3qwgD
D3Kon+28YGWNgz4ootT4QTwQGwUAtZrz+0iTyufQWRvnELBGj7fg6xZ+wEKuaC6VyQZb20IWsJZm
z9ocbAbZlycTo+rXDv2bogmR7d+PmIIovQTyArEV1bQeD/FYVDOpyXdpvKpT2jjrCAZdUNrOaaaa
sMQ+cBJtzQdH+g+zUZ6MLUnZqcGMAu5kIuGX8sbxqEYTWkR3j9mxlOJFoYQyZp1M5ggUSrwgITiZ
CMfIUYKNDTvU6OqYDKPprhdC4igGZYrvVVXpIKx1A2wzVGtsxtppWu7QjpgpCHFTs74VTmGkaHWb
yCJZEQoDF6U2+cmtLKwh8omHA6vnDa/JhRGBAmKciDG+bzaJ/36uH0o2PX2+4qBMm9aw4Dk5JX6v
GA2QFtvyJZX7QUnBMpmRDWzaDcV9RQ9AvDPjkQ+s4Ibm6uYpc36waGiUYWoQEQrYVgfaCvjphReP
YTja54rb35E5h68u4hbXC0fWl/vJpVP3GOC3Db40VwO5Z9pkOwTyA0/BXPQ4+IOxdYV4qryzTt1e
NOb854di69upFwYy7mL8PZcrMo/go5J8r7/KXCWWr/neQtPfd3Y3ie8Qn1o+U2PuV9TB9MKtgh9T
/AuzcnZ24thXraYLgeJ6bWUHvz/lbZGLLMp8Y6E4pk3U7kLgMBdtUJirOCqBpc1kqK9TPFaoNcBW
7JAbJFEzhjn/jOeP6xviC5VHXMCaKrV94aEexv0esBph6nkz5lQMNMwKV8I87kRm9SjFuwRpL+Yo
DcLhrQtv84XHbU/6kV+YwkHJqJLSOfFl7O8e2De+srm1PZzzWeGA5mu+ju6DRwYym+Yqfxv5eYLH
3F2WKS+BoNAH1PYZXH0UC7eCGxSdZocH21NIuyQfamcfNCf5HL5yQlDYodwRqQYx4CvLvvWqliWd
qkInVPfDBnEH/RB6v5MKA2s7iy+8G0dFu/5ZbXtqj4lFjdd2c2oES908ZXJSa58v90/ZBB4eNM3T
PIlJurgdOWASJLkPX+TYo1oRoBGIL8nV26CaJwlKNZDPpxlj+JhGfJBRpgcFAhhYMwQFiGlbbHz0
RpfvJjaqaVJjc8SlNI8GmS71Ptc0Ce9INoXCtaw7ypXNUfMgxTakf0j091taCDV+n9U1cK5LFvbR
eESwljoZMqJGWGQm4yPH4awnL9xSvqwhwJ9I6WtCv/ZQh5ZtcHD3TkGP6Te/anKenrYp5IC08XHL
s2THgMG/QFzEmgiCG7LjTdlnF+xRr/DVees/jBI/OeDieNaeVf4EcayQIBKCzkp1EM0CSwbkxGFh
Onekmf+C+CEIn6+6vKMWvnJm6VHdNPVgnGHjid5wlTRNBx+rQ7DJocc4mZdMPWda3RfEksQ7yk6g
EVnIwHeWouxANmymTXGmo46B5qwjJuCsUE0/Yc/St8egL3I8PoFyiDlx1yhx+I7yNrFV67Yuerb7
M/7Q6Zb0OCCxJLMn0l4t4kVTPeIGl/Zi9d956isymf10EFZkH+9bSidi3vDzn7rguLXcOzP0De+2
/2hgRZOCjcKn7gFg6xWGh+tpr5BdGeKPMvt06WqQKzrpJTRxlL/toBB7shLfITBqoEvwui3RL1bb
qtNhDOEhKdVbWjni/nKhgrC4AoJBv60tTa0SqOZPSs/kI67MmO5kkXiG3boxqMVwfbmqlTcAkw72
0lKPypYVsPydub301lCaVxlWJY7NyALPDCUM9wqPH189qZbBUTQW8JZ1dp+b9Qh/JANGiyPa6EMT
p3iLupKjrNErqYNzTjoeNxIUwH21OfOt2rSfVHZU2YaZrxbrhZmlrBFY+ewLGLt+zDyrrvLQig5y
xKU1xqgn0xEii+Pypn4Bur8IWnCGXiXhJuylEZoxGJZEjyVv8j1h9AQHvwJwaPC9oWsREng1kOC9
dRcjAT6t8xmXhRVhWkYLHsPQOJXJFo3iSJGa1hG6/5Y2xdNApJB0aERnw6HGJdr64JmvlRzV4esv
ljOSSfc6mBq/amvZnOz8WFXupX6yO0D52jxqrhcYdVuvaHW448Euu/lif2PkvwmhPovr7qVLmoLA
lnaayk2LNPebKqye85O+ZlZuM6aYcbFgGs0KX7lQZoIwy1nOYZHo4yujOjOjEUklUW2gUcE2u5Hg
rUngtAulQWBs1lTzH23GOvxuUzDWic5NV72Nlye2Eg7PT6kmQOaYT5vF35ip79bjJ0SqZHCjBK/Z
L7cbI/Xr622YtKJfGNvGvEatwwPLrg3CmhrmXJ0CRCYahBMDqXiUaU1JTx6FS9cWKU5MoIusuZo8
CzGYQu+ukQUKT+ZZ8k7F0HYhh/lR/wi75hKO0yoryKLtjw75Tk2lebajHGyC7AH9C4lkBZpX5iG8
FtVudbgupY/ZXL1hZfIhXxHJA9/AZICOynoVAg2OqXjCoD6Xg+Dx/hoHI+AUlQ5uAdWiDgcTlKDg
Bb2olWHXLlipsOd2Ep8ksbCJD0n8NyYa1HpyGTCzsk/FcC7+0Tkn94w9vFeLCLSXMez9MJhzT+OU
qH4BphIUY8lypVoBUxRmIDBfpcnzldqRMtZUO5itKk1yOINVyx5iKPlpSUpprlxlkajcxAdkDq5F
TQdURQuQDAbUrNAhO2v1EMtJp/5on5/9QSMAq9VIAfKm/gTtB45HU+0grSmGBynichpjgBNgnoiZ
aMBu2vG59AhN8k0NsOIXUOsR0qSHCcxWeGJtqJiGLrqjkLpPmRfYpVu5MpP9wLAacGoc5ngyrUaP
nesUpicJLavqngT+WUUVRQSBcq0JQ0SWjnLCI8N2PykgI5VAcl19TYUElO37ZSiF/WUKNrhKoa6g
0OQf/xFJRr4FQoaYQyodZJojvPEmJird9xS7lb3SfYHmKoW3OYQStvAHtBBXA5IGEEnf16wuHyT0
Vk3RVWMiiUJ+Wj3UcVDRd4xwx9saR6EAVZJJK09neJTu3mXnRBTeOWxO6ZAMG1iZW+ihHS2AGw87
7gd8TZz3irSWL8+OKzcE6+RyMfhr236l/RTVoQ+ejATPY77gFMnXmmHs1MREHPCzZyymdYGUvW21
5F74ULrVZKQMF44tBpkJMkNLYB7OmieSi2NoF9SLiNbPP5mbERZ3St3yVbeEAQ1zyNtxQYtcK3z1
TKH+Qg3BQ9Irh/owD7x2DfRtJtgc0+BHuCcIK4D9160IQ4iPzPgX+A4Iu/rZ/suw55bTMJ0Naiui
muY3ekA5Fe29G3iR3UwKKrG+bR5FPRGIDoQukJe2UPs6jzSypVWlZKybbX25E0cnHw3+kcIUFkbd
JLGmOHePzpW4qK5DdbToCNq/RREujJi6o1CBabs+Vr9DcaFoIAMYVTWE8yoIMO1AE13GkRlBpqCt
Zk/ouAWz4vc4K+V39WhL/eionyh0bwTkHds9lno4P6ZSqIYtTiueOCole1R4t54oxdRvIeg9e0kV
4WfeqJdFsitbM1qBSpvBR4I0KHLE9wqJlR9KXRphQ2CnO5DSv1VEmK/lwTC0tWGcnPvoQiGTrmK4
ivBd2yCtyOUvNzmRRZPkcCJ2wi/WEOzXj/PRW0PXnWu4Z6xzVzXzJ6mkq1VrehX2Z1PlxLWOvakl
O/HRfzuh28Jd85lXd4T9jywlS5KsA7x3rxBiKgVC2KxNIoet9Tf5axXyqEdR8BXTnuh4upq78/CZ
0OXQ+Bwa1DFpVux2VBx/S4RTQCmKwIxEJP2tNm0iCwonfzmUgoefKZaPeUBs9PZMtF/kG9IgszQM
Z4AylRH2yzTDaW1e7N5MoKIWHh8ChQ/elrLqSX+vGYNMHlCxNwCsYJEkBQ8FlOQSTizt/p98yOyB
PsQw0RB3uRcrHs+N5InoXCdBWUluokt6yqeOC+rVLWIa+FrWhf7LFZe9f3E8YxppQqKSPa0i0OEv
7sJdBm0/phGyctWvkyjOkMARW0YqY3Cpe+bGSKsU4jjE6qQ00ufqEGTvnPw5BFZlhLuVQWmbuX08
VIvB6z1DIenEuq3iRmLAiG9JkrKckv33RDyLuNwc6ztEOAp7lvpnQ+/VJJsdNOibC86Yyi44A7GF
JTOnhmmum/EusJRsFu2oBWL0PJ7b9PN3gkx95IhjeWs95f+tCY2ZqM78PNkIFP85YZxzmevwvsFL
1BdQRQVZx5pSP7tuDcDLKEiEaMdfUkpW5BYoagzJqqX0j1addpZewrHUFyeko5d3layfszEhf31J
/3FLR3eSSaNu3n2bnPldfbWZ/SgvOVGMkfE9hABylYbCgBoM2PslD693JNPRtemxeaHm76+fixFv
8MTYV85V3IEiHlsE/crCChw4PiK4Uu5CYkzEFdx3JWhzngwgxbuxddqV18xhrV+kRghQ/yB2kEsk
L4r7itTCICZ9SM5irK0wpa+X1dYFgrMgdxLyaxV5jguzLt02sHGJl2QYZo7e0JYt01Nb9V/cRByj
+JIFp2m5Or9U62bIhHTHmsZWruLDH6ypj0fo3zHHM8VkQJEFq2aD7tJsB+l5tdjgQzREJTJGgU/O
DMzmGq8xsJzJRkxgq+dnSizoVbD2DZ30y2W32eGCVh6OKz/0gCBdAabZuo7dTpt7rGpMfPBqeb0D
wDJCR6Q7NmQIt/AVOQyi0Y0jxglyrsV5HqVlZ1irGBC6IuDjHzVnlAVHRQ8YP2o7t/kKGtubhS+Q
IKXpO5QN4KU6iPcGi24lhTh6zcfoj+ApVDrVau1RHrmndqS7KJOqteN6GTzdD0rkBiFJc12Sa/fV
ToMn0tx+GdvDfXLID1TpaHZyu6iDz7Tu0RKV8MJtoDj1yZjnCCF0uoaLwb4bfo5AKaNypT8iA0yv
/YsnrvOM9j1Q90vKDR3NXlviZd6GXZsWNM7oKEsGW4bEIHHubufyrEOUb1hyOrFDzDdl9DjIuCGJ
SNEx/GKxhe3GnXFhWNaGdIwlUkAwIKDgdaBr5ytdH2OcPyjPfzSlIq9I+bKh8ePM9S1hablyJssZ
9p1+BYnEnqow1N4m+1yR+khf3OiiMSNhvG2FjA/RUGuHHj1mQVJ6BCeAFkKltPUnMJvYq4A5JMqq
CM9wcu9Z0otI6ZmQNPi+vuB7HUP5f1fCnVt0tLyIA4uX4Cs/PCWCmoNXdkZf8Jjy0JV2Lh8zLTpR
jY8uw0ksIz5tlZ+e82y7imPLYukkvsz+AbdjdcSAyMn7bvnSGR0Z3+QRgi932mZDFxvSIqrPHi/L
xwhHW0nrDPMlPU1sdfHlK3qjXnRHFNhkdfCzJyshOoqhZKao83TN8XLan4WLt1FJjoZDGP+CAuFj
dpTdrhPNWGMsgBqZDiN4GKxd+PeA1gYQlT+ls0VW7jFZnL87HjHl+IjH9GBmCKnBFbc0KABi2kkJ
YRTFI3SXswxWn5JF8oXiOgItm2I3Zewdox4R26586djr3EV4QR2N7GOFnfErPH8lMSBsapOeJ07r
k5LlKQ9raPx1Rlblg18GuHwDbphoEfR/Y6UV6rVLg1JWG2f0zVF+uE+/apNqpXW5Ldl8cqF8k1Nb
louAyIgc2gfe1UENBWpKwPuOggQ2glxWjba2sWTndirxyPxHTlf0bLha7fPFD+8TQ91qDxTHzdkH
iK2QKld5xLt5abgPHMiAM5wGnCWg0xqqKL+GsaAH6JxgESEyxeA5CjfBtMBA886wsFcF5iPZvPsc
s8UoFBllR/wdUprzVw8hD7SWlAF43xLG2ZTvVyFLfQHAmC8GYAEugbZk9kcghGzKCYEzme6oVB2G
7hLyNhFePKN1/ZaGeZBloPW8PrPf3xYUXT821YCfDpOE9+WN2S8O/DHPxKmAgv74jOUnP4kF7+g8
ebfuDxNOqJ4Mk6OXKOsWDMu3/7sr9mpBvdOcH/kR2cygZ3BjZbZOO98XVJmiwvBBqOMfBdkklkGT
aJ4hw+YTmgddWC8nWEHTC/oMXGH3PS5rZe4RRpR74FDm90+nT/TllGUjqbHyIswKcGIFait03awx
v8xwiQBt7JhbRu0Cuce4UMCJW0nZDDtQBH8zUgnfmF/rkik792dL9q54Hshl72JtV7dLdI39ws3x
d1US2HFFXB6m9a5FoO2DYRxM/mAut/BzzxazXq8cPZ3PbfFxi4qYxIyItwVVw0j12CfpWM7ungDF
WQMTfCtbClif0rDEeLsx9fXB4CRs80wOeaAGYR1gedj8WXJcM6lJDcqjHyGF0EO/NG4cSrzszGaw
+PR9SAqMZrik1kRj+OTxq9TXjh3dM5WcsM1lE6sxmtXTohVzM017uouCJAt9cpc9t23XRkwPzJd8
u3sdTrRHgeYrl+w1hjrOHsUFd7/EZVOImXbB3xAXN7KtXepr6T3WGNC3JtCXE/6NofY7fpbBGS6E
IN24qpBfUEB09zdrrF0jvCuLUIyr2wtr1CEVCsH5lmblnIaj+y6zpnvAPecoFpPkCDBPpTUOIi+D
G/FqLNlwT3gC/nRhKnowI8uXO2wzG0Vcwz3TeNkJLz0W4/kbkd9WMsPjnyE03uyi1uNE8KXkyl4K
8DdleZNeg7Lj9ADIPJsv3HdxK1QwM/2KTQ1o45eUxLe6wBTX9AURTwV6lnUNNFA636Nwz+FTYU0v
r80yZOcxcR/8x5dEajux7s2iMRnZzepR2bCNsOMWGB6dov2gIahDFNj8VgMKPwuN8jIls32DABbx
hi3qq6InoWlsPLzU1kID91ovLvytafc+9MTn6MGrEE1cNxqGtPKg3lfwjlZLnsqRPbArZn4deV0x
eK+7B5dfz7hhgArQaQQXhKCGjY2Z/TEo1LIf9UjxmyknynVeyPbx9XR65aRbUxIuWb5n5UsUUZU+
KoGFHgm52/3Ok2Y+6WKCXtLnCSvx66Bh8kjGmRRRFlfzjPugzsdoxCaAWjrWxP9+BvMay7OwDXiQ
Hokn7omSYWV0VwIZpWhgFxES3kv1NWTG/i0rK7/pC49cFAkFO2bBJWu3ARW2nMI2wlVnwR2q0CR6
jitdjeDBRK7tfcivdkZqC4g5jT0ewAuz7b50NpaX73DVn17TBZxIEH+8t1PTcb7WqOTOnuB7TqgF
PN6WO9AaHLhf9otgAIBcdhzKci5mPMNXv153aidP81rPEWK+wt1whSTM3gnTIZqg/ZzJQHGjJ3/V
a00MHVbehcG29viSic8ysVDO6pdvpC4FbXztK7oBNHeLX9ZAZC6mNMBNEymbnoPY2BZhCi/3ghJu
PmiiGCOSakzfaAXUPppYamykDJxtUhA8Aj8VEvGQcy15yiA50Wq8NCR3XqkMr7Jfws8lOgKGvXjX
vWZt+U9Fvyn31vsdtd4TiIcVdFwTc3NK0kMCsb3X0Y/GjrhiREfuuvzpu2SqaaiPaVxJ79jsNJTN
Hr+aI83Srj6vZIy+geNXtpEXvqrx3ZelpKCnR8sem6kgk3k/LuNYJmu2xw/OvebHjq3w5dSae6jp
E3DfcTYhP8fooYyEyPukQrRqTD1vFvPTQsUO2hzRAKPR3aPhk49H3AxGie75g7qTQrASZXD/DaBU
yqBTfRcfES2AUnj1i8QPxxDT32omox9PY+BZlhR8/tOJTxJtX9A+NEp/mueCM4Ux6+jKTgIFCgVU
xq+FJ0F6FLGWrBVYrIEsD37fx5IsRncq0+7HHtIaxKk3pLToYxSCxd1ERsL5Vk3n7nqn2loO0LJy
68hFHbeEUKAu6yO4mD7MUG9OYWi/gHsmTK4/dWRyTc3en4CzgY4vjJ1ckNA8N0T5hYqTdzwDJr2I
EosU4n5rUk1zB8FJVdF4oq9OT7VupEWcfJoLNS7sDMCdnQh/roPQ06x1Xn6c2gAygCv3vJGHHl1+
r8UXwD0cYkeyDTlzm3FxH5DStOX5OP5WgTlPWzG8TA9WiqEDroS5lWfkAoT0EhyimzVlurQj0NXP
vl5CNa+TO6x8a9oppuAhimV7yGhEBBCuAaGUBW3nwl/kJ08hWCaXvUirbg==
`protect end_protected
