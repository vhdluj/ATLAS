------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gtx_quad_no_buffer_exdes.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gtx_quad_no_buffer_exdes
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity gtx_quad_no_buffer_exdes is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;    -- specifies lane with unique start frame ch
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;  -- specifies amount of data in BRAM
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";    -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 1;             -- Set to 1 for simulation
    STABLE_CLOCK_PERIOD                     : integer   := 16; 
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets
);
port
(
    Q0_CLK1_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_PAD_P_IN               : in   std_logic;
    DRP_CLK_IN                              : in   std_logic;
    TRACK_DATA_OUT                          : out  std_logic;
    RXN_IN                                  : in   std_logic_vector(3 downto 0);
    RXP_IN                                  : in   std_logic_vector(3 downto 0);
    TXN_OUT                                 : out  std_logic_vector(3 downto 0);
    TXP_OUT                                 : out  std_logic_vector(3 downto 0)
    
);


end gtx_quad_no_buffer_exdes;
    
architecture RTL of gtx_quad_no_buffer_exdes is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gtx_quad_no_buffer,gtwizard_v2_6,{protocol_file=Start_from_scratch}";

--**************************Component Declarations*****************************


component gtx_quad_no_buffer_init
generic
(
    -- Simulation attributes
    EXAMPLE_SIM_GTRESET_SPEEDUP    : string    := "FALSE";    -- Set to 1 to speed up sim reset
    EXAMPLE_SIMULATION             : integer   := 0;          -- Set to 1 for simulation
    STABLE_CLOCK_PERIOD            : integer   := 16; 
    EXAMPLE_USE_CHIPSCOPE          : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT0_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_RX_MMCM_RESET_OUT                   : out  std_logic;

    --_________________________________________________________________________
        --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt0_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt0_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt0_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt0_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt0_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gtxrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    gt0_rxpmareset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt0_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt0_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gtxtxn_out                          : out  std_logic;
    gt0_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
   
    --_________________________________________________________________________
        --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt1_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt1_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt1_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt1_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt1_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gtxrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    gt1_rxpmareset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt1_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt1_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt1_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gtxtxn_out                          : out  std_logic;
    gt1_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
   
    --_________________________________________________________________________
        --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt2_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt2_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt2_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt2_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt2_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gtxrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    gt2_rxpmareset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt2_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt2_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt2_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gtxtxn_out                          : out  std_logic;
    gt2_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
   
    --_________________________________________________________________________
        --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt3_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt3_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt3_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt3_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    gt3_gtxrxp_in                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gtxrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    gt3_rxpmareset_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt3_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt3_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt3_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gtxtxn_out                          : out  std_logic;
    gt3_gtxtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
   

    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    gt0_gtrefclk0_common_in                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    gt0_qplllock_out                        : out  std_logic;
    gt0_qplllockdetclk_in                   : in   std_logic;
    gt0_qpllpd_in                           : in   std_logic;
    gt0_qpllreset_in                        : in   std_logic


);
end component;

component gtx_quad_no_buffer_GT_USRCLK_SOURCE 
port
(
    Q0_CLK1_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_OUT                    : out  std_logic;
 
    GT0_TXUSRCLK_OUT             : out std_logic;
    GT0_TXUSRCLK2_OUT            : out std_logic;
    GT0_TXOUTCLK_IN              : in  std_logic;
    GT0_TXCLK_LOCK_OUT           : out std_logic;
    GT0_TX_MMCM_RESET_IN         : in std_logic;
    GT0_RXUSRCLK_OUT             : out std_logic;
    GT0_RXUSRCLK2_OUT            : out std_logic;
    GT0_RXOUTCLK_IN              : in  std_logic;
    GT0_RXCLK_LOCK_OUT           : out std_logic;
    GT0_RX_MMCM_RESET_IN         : in std_logic;
 
    GT1_TXUSRCLK_OUT             : out std_logic;
    GT1_TXUSRCLK2_OUT            : out std_logic;
    GT1_TXOUTCLK_IN              : in  std_logic;
    GT1_TXCLK_LOCK_OUT           : out std_logic;
    GT1_TX_MMCM_RESET_IN         : in std_logic;
    GT1_RXUSRCLK_OUT             : out std_logic;
    GT1_RXUSRCLK2_OUT            : out std_logic;
    GT1_RXOUTCLK_IN              : in  std_logic;
    GT1_RXCLK_LOCK_OUT           : out std_logic;
    GT1_RX_MMCM_RESET_IN         : in std_logic;
 
    GT2_TXUSRCLK_OUT             : out std_logic;
    GT2_TXUSRCLK2_OUT            : out std_logic;
    GT2_TXOUTCLK_IN              : in  std_logic;
    GT2_TXCLK_LOCK_OUT           : out std_logic;
    GT2_TX_MMCM_RESET_IN         : in std_logic;
    GT2_RXUSRCLK_OUT             : out std_logic;
    GT2_RXUSRCLK2_OUT            : out std_logic;
    GT2_RXOUTCLK_IN              : in  std_logic;
    GT2_RXCLK_LOCK_OUT           : out std_logic;
    GT2_RX_MMCM_RESET_IN         : in std_logic;
 
    GT3_TXUSRCLK_OUT             : out std_logic;
    GT3_TXUSRCLK2_OUT            : out std_logic;
    GT3_TXOUTCLK_IN              : in  std_logic;
    GT3_TXCLK_LOCK_OUT           : out std_logic;
    GT3_TX_MMCM_RESET_IN         : in std_logic;
    GT3_RXUSRCLK_OUT             : out std_logic;
    GT3_RXUSRCLK2_OUT            : out std_logic;
    GT3_RXOUTCLK_IN              : in  std_logic;
    GT3_RXCLK_LOCK_OUT           : out std_logic;
    GT3_RX_MMCM_RESET_IN         : in std_logic;
    DRPCLK_IN                          : in  std_logic;
    DRPCLK_OUT                         : out std_logic
);
end component;




component gtx_quad_no_buffer_GT_FRAME_GEN 
generic
(
     WORDS_IN_BRAM    : integer := 512
);
port
(
    -- User Interface
    TX_DATA_OUT             : out   std_logic_vector(79 downto 0);
    TXCTRL_OUT              : out   std_logic_vector(7 downto 0); 
    -- System Interface
    USER_CLK                : in    std_logic;      
    SYSTEM_RESET            : in    std_logic
); 
end component;

component gtx_quad_no_buffer_GT_FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    RXCTRL_WIDTH             : integer := 2; 
    WORDS_IN_BRAM            : integer := 256;
    CHANBOND_SEQ_LEN         : integer := 1;
    COMMA_DOUBLE             : std_logic_vector(15 downto 0) := x"f628";
    START_OF_PACKET_CHAR     : std_logic_vector(31 downto 0) := x"060504bc"
);
port
(
    -- User Interface
    RX_DATA_IN               : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    RXCTRL_IN                : in  std_logic_vector((RXCTRL_WIDTH-1) downto 0); 
    RXENMCOMMADET_OUT        : out std_logic;
    RXENPCOMMADET_OUT        : out std_logic;
    RX_ENCHAN_SYNC_OUT       : out std_logic;
    RX_CHANBOND_SEQ_IN       : in  std_logic;

    -- Control Interface
    INC_IN                   : in  std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCHB_OUT       : out std_logic;
    RESET_ON_ERROR_IN        : in  std_logic;


    -- Error Monitoring
    ERROR_COUNT_OUT          : out std_logic_vector(7 downto 0);

    -- Track Data
    TRACK_DATA_OUT           : out std_logic;

 

    -- System Interface
    USER_CLK                 : in std_logic;       
    SYSTEM_RESET             : in std_logic
);
end component;

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

    signal   gt0_txfsmresetdone_i            : std_logic;
signal   gt0_rxfsmresetdone_i            : std_logic;
    signal   gt0_txfsmresetdone_r            : std_logic;
    signal   gt0_txfsmresetdone_r2           : std_logic;
signal   gt0_rxresetdone_r               : std_logic;
signal   gt0_rxresetdone_r2              : std_logic;
signal   gt0_rxresetdone_r3              : std_logic;


    signal   gt1_txfsmresetdone_i            : std_logic;
signal   gt1_rxfsmresetdone_i            : std_logic;
    signal   gt1_txfsmresetdone_r            : std_logic;
    signal   gt1_txfsmresetdone_r2           : std_logic;
signal   gt1_rxresetdone_r               : std_logic;
signal   gt1_rxresetdone_r2              : std_logic;
signal   gt1_rxresetdone_r3              : std_logic;


    signal   gt2_txfsmresetdone_i            : std_logic;
signal   gt2_rxfsmresetdone_i            : std_logic;
    signal   gt2_txfsmresetdone_r            : std_logic;
    signal   gt2_txfsmresetdone_r2           : std_logic;
signal   gt2_rxresetdone_r               : std_logic;
signal   gt2_rxresetdone_r2              : std_logic;
signal   gt2_rxresetdone_r3              : std_logic;


    signal   gt3_txfsmresetdone_i            : std_logic;
signal   gt3_rxfsmresetdone_i            : std_logic;
    signal   gt3_txfsmresetdone_r            : std_logic;
    signal   gt3_txfsmresetdone_r2           : std_logic;
signal   gt3_rxresetdone_r               : std_logic;
signal   gt3_rxresetdone_r2              : std_logic;
signal   gt3_rxresetdone_r3              : std_logic;


signal   reset_pulse                     : std_logic_vector(3 downto 0);
    signal   reset_counter  :   unsigned(5 downto 0) := "000000";


--**************************** Wire Declarations ******************************
    -------------------------- GT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GT0  (X0Y0)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt0_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt0_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpen_i                     : std_logic;
    signal  gt0_drprdy_i                    : std_logic;
    signal  gt0_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt0_loopback_i                  : std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    signal  gt0_rxpd_i                      : std_logic_vector(1 downto 0);
    signal  gt0_txpd_i                      : std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt0_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt0_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt0_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt0_rxdata_i                    : std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt0_rxdisperr_i                 : std_logic_vector(3 downto 0);
    signal  gt0_rxnotintable_i              : std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    signal  gt0_gtxrxp_i                    : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt0_gtxrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt0_rxdlyen_i                   : std_logic;
    signal  gt0_rxdlysreset_i               : std_logic;
    signal  gt0_rxdlysresetdone_i           : std_logic;
    signal  gt0_rxphalign_i                 : std_logic;
    signal  gt0_rxphaligndone_i             : std_logic;
    signal  gt0_rxphalignen_i               : std_logic;
    signal  gt0_rxphdlyreset_i              : std_logic;
    signal  gt0_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt0_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt0_rxmcommaalignen_i           : std_logic;
    signal  gt0_rxpcommaalignen_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt0_rxlpmhfhold_i               : std_logic;
    signal  gt0_rxlpmlfhold_i               : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt0_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt0_gtrxreset_i                 : std_logic;
    signal  gt0_rxpmareset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt0_rxcharisk_i                 : std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt0_rxresetdone_i               : std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    signal  gt0_txpostcursor_i              : std_logic_vector(4 downto 0);
    signal  gt0_txprecursor_i               : std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt0_gttxreset_i                 : std_logic;
    signal  gt0_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt0_txdlyen_i                   : std_logic;
    signal  gt0_txdlysreset_i               : std_logic;
    signal  gt0_txdlysresetdone_i           : std_logic;
    signal  gt0_txphalign_i                 : std_logic;
    signal  gt0_txphaligndone_i             : std_logic;
    signal  gt0_txphalignen_i               : std_logic;
    signal  gt0_txphdlyreset_i              : std_logic;
    signal  gt0_txphinit_i                  : std_logic;
    signal  gt0_txphinitdone_i              : std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    signal  gt0_txdiffctrl_i                : std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt0_txdata_i                    : std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt0_gtxtxn_i                    : std_logic;
    signal  gt0_gtxtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt0_txoutclk_i                  : std_logic;
    signal  gt0_txoutclkfabric_i            : std_logic;
    signal  gt0_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt0_txcharisk_i                 : std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt0_txresetdone_i               : std_logic;

    --________________________________________________________________________
    --________________________________________________________________________
    --GT1  (X0Y1)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt1_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt1_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt1_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt1_drpen_i                     : std_logic;
    signal  gt1_drprdy_i                    : std_logic;
    signal  gt1_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt1_loopback_i                  : std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    signal  gt1_rxpd_i                      : std_logic_vector(1 downto 0);
    signal  gt1_txpd_i                      : std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt1_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt1_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt1_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt1_rxdata_i                    : std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt1_rxdisperr_i                 : std_logic_vector(3 downto 0);
    signal  gt1_rxnotintable_i              : std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    signal  gt1_gtxrxp_i                    : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt1_gtxrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt1_rxdlyen_i                   : std_logic;
    signal  gt1_rxdlysreset_i               : std_logic;
    signal  gt1_rxdlysresetdone_i           : std_logic;
    signal  gt1_rxphalign_i                 : std_logic;
    signal  gt1_rxphaligndone_i             : std_logic;
    signal  gt1_rxphalignen_i               : std_logic;
    signal  gt1_rxphdlyreset_i              : std_logic;
    signal  gt1_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt1_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt1_rxmcommaalignen_i           : std_logic;
    signal  gt1_rxpcommaalignen_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt1_rxlpmhfhold_i               : std_logic;
    signal  gt1_rxlpmlfhold_i               : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt1_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt1_gtrxreset_i                 : std_logic;
    signal  gt1_rxpmareset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt1_rxcharisk_i                 : std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt1_rxresetdone_i               : std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    signal  gt1_txpostcursor_i              : std_logic_vector(4 downto 0);
    signal  gt1_txprecursor_i               : std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt1_gttxreset_i                 : std_logic;
    signal  gt1_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt1_txdlyen_i                   : std_logic;
    signal  gt1_txdlysreset_i               : std_logic;
    signal  gt1_txdlysresetdone_i           : std_logic;
    signal  gt1_txphalign_i                 : std_logic;
    signal  gt1_txphaligndone_i             : std_logic;
    signal  gt1_txphalignen_i               : std_logic;
    signal  gt1_txphdlyreset_i              : std_logic;
    signal  gt1_txphinit_i                  : std_logic;
    signal  gt1_txphinitdone_i              : std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    signal  gt1_txdiffctrl_i                : std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt1_txdata_i                    : std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt1_gtxtxn_i                    : std_logic;
    signal  gt1_gtxtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt1_txoutclk_i                  : std_logic;
    signal  gt1_txoutclkfabric_i            : std_logic;
    signal  gt1_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt1_txcharisk_i                 : std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt1_txresetdone_i               : std_logic;

    --________________________________________________________________________
    --________________________________________________________________________
    --GT2  (X0Y2)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt2_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt2_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt2_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt2_drpen_i                     : std_logic;
    signal  gt2_drprdy_i                    : std_logic;
    signal  gt2_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt2_loopback_i                  : std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    signal  gt2_rxpd_i                      : std_logic_vector(1 downto 0);
    signal  gt2_txpd_i                      : std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt2_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt2_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt2_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt2_rxdata_i                    : std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt2_rxdisperr_i                 : std_logic_vector(3 downto 0);
    signal  gt2_rxnotintable_i              : std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    signal  gt2_gtxrxp_i                    : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt2_gtxrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt2_rxdlyen_i                   : std_logic;
    signal  gt2_rxdlysreset_i               : std_logic;
    signal  gt2_rxdlysresetdone_i           : std_logic;
    signal  gt2_rxphalign_i                 : std_logic;
    signal  gt2_rxphaligndone_i             : std_logic;
    signal  gt2_rxphalignen_i               : std_logic;
    signal  gt2_rxphdlyreset_i              : std_logic;
    signal  gt2_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt2_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt2_rxmcommaalignen_i           : std_logic;
    signal  gt2_rxpcommaalignen_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt2_rxlpmhfhold_i               : std_logic;
    signal  gt2_rxlpmlfhold_i               : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt2_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt2_gtrxreset_i                 : std_logic;
    signal  gt2_rxpmareset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt2_rxcharisk_i                 : std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt2_rxresetdone_i               : std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    signal  gt2_txpostcursor_i              : std_logic_vector(4 downto 0);
    signal  gt2_txprecursor_i               : std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt2_gttxreset_i                 : std_logic;
    signal  gt2_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt2_txdlyen_i                   : std_logic;
    signal  gt2_txdlysreset_i               : std_logic;
    signal  gt2_txdlysresetdone_i           : std_logic;
    signal  gt2_txphalign_i                 : std_logic;
    signal  gt2_txphaligndone_i             : std_logic;
    signal  gt2_txphalignen_i               : std_logic;
    signal  gt2_txphdlyreset_i              : std_logic;
    signal  gt2_txphinit_i                  : std_logic;
    signal  gt2_txphinitdone_i              : std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    signal  gt2_txdiffctrl_i                : std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt2_txdata_i                    : std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt2_gtxtxn_i                    : std_logic;
    signal  gt2_gtxtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt2_txoutclk_i                  : std_logic;
    signal  gt2_txoutclkfabric_i            : std_logic;
    signal  gt2_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt2_txcharisk_i                 : std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt2_txresetdone_i               : std_logic;

    --________________________________________________________________________
    --________________________________________________________________________
    --GT3  (X0Y3)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt3_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt3_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt3_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt3_drpen_i                     : std_logic;
    signal  gt3_drprdy_i                    : std_logic;
    signal  gt3_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt3_loopback_i                  : std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    signal  gt3_rxpd_i                      : std_logic_vector(1 downto 0);
    signal  gt3_txpd_i                      : std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt3_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt3_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt3_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt3_rxdata_i                    : std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt3_rxdisperr_i                 : std_logic_vector(3 downto 0);
    signal  gt3_rxnotintable_i              : std_logic_vector(3 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    signal  gt3_gtxrxp_i                    : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt3_gtxrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt3_rxdlyen_i                   : std_logic;
    signal  gt3_rxdlysreset_i               : std_logic;
    signal  gt3_rxdlysresetdone_i           : std_logic;
    signal  gt3_rxphalign_i                 : std_logic;
    signal  gt3_rxphaligndone_i             : std_logic;
    signal  gt3_rxphalignen_i               : std_logic;
    signal  gt3_rxphdlyreset_i              : std_logic;
    signal  gt3_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt3_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt3_rxmcommaalignen_i           : std_logic;
    signal  gt3_rxpcommaalignen_i           : std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt3_rxlpmhfhold_i               : std_logic;
    signal  gt3_rxlpmlfhold_i               : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt3_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt3_gtrxreset_i                 : std_logic;
    signal  gt3_rxpmareset_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt3_rxcharisk_i                 : std_logic_vector(3 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt3_rxresetdone_i               : std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    signal  gt3_txpostcursor_i              : std_logic_vector(4 downto 0);
    signal  gt3_txprecursor_i               : std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt3_gttxreset_i                 : std_logic;
    signal  gt3_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt3_txdlyen_i                   : std_logic;
    signal  gt3_txdlysreset_i               : std_logic;
    signal  gt3_txdlysresetdone_i           : std_logic;
    signal  gt3_txphalign_i                 : std_logic;
    signal  gt3_txphaligndone_i             : std_logic;
    signal  gt3_txphalignen_i               : std_logic;
    signal  gt3_txphdlyreset_i              : std_logic;
    signal  gt3_txphinit_i                  : std_logic;
    signal  gt3_txphinitdone_i              : std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    signal  gt3_txdiffctrl_i                : std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt3_txdata_i                    : std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt3_gtxtxn_i                    : std_logic;
    signal  gt3_gtxtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt3_txoutclk_i                  : std_logic;
    signal  gt3_txoutclkfabric_i            : std_logic;
    signal  gt3_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt3_txcharisk_i                 : std_logic_vector(3 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt3_txresetdone_i               : std_logic;

    --____________________________COMMON PORTS________________________________
    ------------------------- Common Block - QPLL Ports ------------------------
    signal  gt0_qplllock_i                  : std_logic;
    signal  gt0_qpllpd_i                    : std_logic;
    signal  gt0_qpllrefclklost_i            : std_logic;
    signal  gt0_qpllreset_i                 : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  gt0_tx_system_reset_c           : std_logic;
    signal  gt0_rx_system_reset_c           : std_logic;
    signal  gt1_tx_system_reset_c           : std_logic;
    signal  gt1_rx_system_reset_c           : std_logic;
    signal  gt2_tx_system_reset_c           : std_logic;
    signal  gt2_rx_system_reset_c           : std_logic;
    signal  gt3_tx_system_reset_c           : std_logic;
    signal  gt3_rx_system_reset_c           : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drpclk_in_i                     : std_logic;
    signal  GTTXRESET_IN                    : std_logic;
    signal  GTRXRESET_IN                    : std_logic;
    signal  QPLLRESET_IN                    : std_logic;

    attribute keep: string;
   ------------------------------- User Clocks ---------------------------------
    signal    gt0_txusrclk_i                  : std_logic; 
    signal    gt0_txusrclk2_i                 : std_logic; 
    signal    gt0_rxusrclk_i                  : std_logic; 
    signal    gt0_rxusrclk2_i                 : std_logic; 
    attribute keep of gt0_txusrclk_i : signal is "true";
    attribute keep of gt0_txusrclk2_i : signal is "true";
    attribute keep of gt0_rxusrclk_i : signal is "true";
    attribute keep of gt0_rxusrclk2_i : signal is "true";
    signal    gt1_txusrclk_i                  : std_logic; 
    signal    gt1_txusrclk2_i                 : std_logic; 
    signal    gt1_rxusrclk_i                  : std_logic; 
    signal    gt1_rxusrclk2_i                 : std_logic; 
    attribute keep of gt1_txusrclk_i : signal is "true";
    attribute keep of gt1_txusrclk2_i : signal is "true";
    attribute keep of gt1_rxusrclk_i : signal is "true";
    attribute keep of gt1_rxusrclk2_i : signal is "true";
    signal    gt2_txusrclk_i                  : std_logic; 
    signal    gt2_txusrclk2_i                 : std_logic; 
    signal    gt2_rxusrclk_i                  : std_logic; 
    signal    gt2_rxusrclk2_i                 : std_logic; 
    attribute keep of gt2_txusrclk_i : signal is "true";
    attribute keep of gt2_txusrclk2_i : signal is "true";
    attribute keep of gt2_rxusrclk_i : signal is "true";
    attribute keep of gt2_rxusrclk2_i : signal is "true";
    signal    gt3_txusrclk_i                  : std_logic; 
    signal    gt3_txusrclk2_i                 : std_logic; 
    signal    gt3_rxusrclk_i                  : std_logic; 
    signal    gt3_rxusrclk2_i                 : std_logic; 
    attribute keep of gt3_txusrclk_i : signal is "true";
    attribute keep of gt3_txusrclk2_i : signal is "true";
    attribute keep of gt3_rxusrclk_i : signal is "true";
    attribute keep of gt3_rxusrclk2_i : signal is "true";
    signal    gt0_txmmcm_lock_i               : std_logic;
    signal    gt0_txmmcm_reset_i              : std_logic;
    signal    gt0_rxmmcm_lock_i               : std_logic; 
    signal    gt0_rxmmcm_reset_i              : std_logic;
    signal    gt1_txmmcm_lock_i               : std_logic;
    signal    gt1_txmmcm_reset_i              : std_logic;
    signal    gt1_rxmmcm_lock_i               : std_logic; 
    signal    gt1_rxmmcm_reset_i              : std_logic;
    signal    gt2_txmmcm_lock_i               : std_logic;
    signal    gt2_txmmcm_reset_i              : std_logic;
    signal    gt2_rxmmcm_lock_i               : std_logic; 
    signal    gt2_rxmmcm_reset_i              : std_logic;
    signal    gt3_txmmcm_lock_i               : std_logic;
    signal    gt3_txmmcm_reset_i              : std_logic;
    signal    gt3_rxmmcm_lock_i               : std_logic; 
    signal    gt3_rxmmcm_reset_i              : std_logic;
    ----------------------------- Reference Clocks ----------------------------
    
signal    q0_clk1_refclk_i                : std_logic;


    ----------------------- Frame check/gen Module Signals --------------------
signal    gt0_matchn_i                    : std_logic;
    
signal    gt0_txcharisk_float_i           : std_logic_vector(3 downto 0);
    
signal    gt0_txdata_float16_i            : std_logic_vector(15 downto 0);
signal    gt0_txdata_float_i              : std_logic_vector(31 downto 0);
    
signal    gt0_track_data_i                : std_logic;
signal    gt0_block_sync_i                : std_logic;
signal    gt0_error_count_i               : std_logic_vector(7 downto 0);
signal    gt0_frame_check_reset_i         : std_logic;
signal    gt0_inc_in_i                    : std_logic;
signal    gt0_inc_out_i                   : std_logic;
signal    gt0_unscrambled_data_i          : std_logic_vector(31 downto 0);

signal    gt1_matchn_i                    : std_logic;
    
signal    gt1_txcharisk_float_i           : std_logic_vector(3 downto 0);
    
signal    gt1_txdata_float16_i            : std_logic_vector(15 downto 0);
signal    gt1_txdata_float_i              : std_logic_vector(31 downto 0);
    
signal    gt1_track_data_i                : std_logic;
signal    gt1_block_sync_i                : std_logic;
signal    gt1_error_count_i               : std_logic_vector(7 downto 0);
signal    gt1_frame_check_reset_i         : std_logic;
signal    gt1_inc_in_i                    : std_logic;
signal    gt1_inc_out_i                   : std_logic;
signal    gt1_unscrambled_data_i          : std_logic_vector(31 downto 0);

signal    gt2_matchn_i                    : std_logic;
    
signal    gt2_txcharisk_float_i           : std_logic_vector(3 downto 0);
    
signal    gt2_txdata_float16_i            : std_logic_vector(15 downto 0);
signal    gt2_txdata_float_i              : std_logic_vector(31 downto 0);
    
signal    gt2_track_data_i                : std_logic;
signal    gt2_block_sync_i                : std_logic;
signal    gt2_error_count_i               : std_logic_vector(7 downto 0);
signal    gt2_frame_check_reset_i         : std_logic;
signal    gt2_inc_in_i                    : std_logic;
signal    gt2_inc_out_i                   : std_logic;
signal    gt2_unscrambled_data_i          : std_logic_vector(31 downto 0);

signal    gt3_matchn_i                    : std_logic;
    
signal    gt3_txcharisk_float_i           : std_logic_vector(3 downto 0);
    
signal    gt3_txdata_float16_i            : std_logic_vector(15 downto 0);
signal    gt3_txdata_float_i              : std_logic_vector(31 downto 0);
    
signal    gt3_track_data_i                : std_logic;
signal    gt3_block_sync_i                : std_logic;
signal    gt3_error_count_i               : std_logic_vector(7 downto 0);
signal    gt3_frame_check_reset_i         : std_logic;
signal    gt3_inc_in_i                    : std_logic;
signal    gt3_inc_out_i                   : std_logic;
signal    gt3_unscrambled_data_i          : std_logic_vector(31 downto 0);

signal    reset_on_data_error_i           : std_logic;
signal    track_data_out_i                : std_logic;
  

    ----------------------- Debug Signals ---------------------------------

    signal  tx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  ila_control_i                   : std_logic_vector(35 downto 0);
    signal  channel_drp_vio_control_i       : std_logic_vector(35 downto 0);
    signal  common_drp_vio_control_i        : std_logic_vector(35 downto 0);
    signal  tx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  tx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);
    signal  ila_in_i                        : std_logic_vector(163 downto 0);
    signal  channel_drp_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  common_drp_vio_async_in_i       : std_logic_vector(31 downto 0);
    signal  common_drp_vio_sync_in_i        : std_logic_vector(31 downto 0);
    signal  common_drp_vio_async_out_i      : std_logic_vector(31 downto 0);
    signal  common_drp_vio_sync_out_i       : std_logic_vector(31 downto 0);

    signal  gt0_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt0_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt0_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);

    signal  gt1_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt1_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt1_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt1_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt1_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt1_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt1_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt1_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt1_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);

    signal  gt2_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt2_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt2_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt2_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt2_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt2_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt2_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt2_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt2_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);

    signal  gt3_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt3_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt3_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt3_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt3_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt3_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt3_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt3_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt3_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);


signal    gttxreset_i                     : std_logic;
signal    gtrxreset_i                     : std_logic;
signal    mux_sel_i                       : std_logic_vector(1 downto 0);

signal    user_tx_reset_i                 : std_logic;
signal    user_rx_reset_i                 : std_logic;
signal    tx_vio_clk_i                    : std_logic;
signal    tx_vio_clk_mux_out_i            : std_logic;    
signal    rx_vio_ila_clk_i                : std_logic;
signal    rx_vio_ila_clk_mux_out_i        : std_logic;    

signal    qpllreset_i                     : std_logic;
    


   function and_reduce(arg: std_logic_vector) return std_logic is
	variable result: std_logic;
    begin
	result := '1';
	for i in arg'range loop
	    result := result and arg(i);
	end loop;
        return result;
    end;


--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
tied_to_ground_i                             <= '0';
tied_to_ground_vec_i                         <= x"0000000000000000";
tied_to_vcc_i                                <= '1';
tied_to_vcc_vec_i                            <= "11111111";

    
  
    
  
    
  
    
  
    gt_usrclk_source : gtx_quad_no_buffer_GT_USRCLK_SOURCE
    port map
   (
        Q0_CLK1_GTREFCLK_PAD_N_IN       =>      Q0_CLK1_GTREFCLK_PAD_N_IN,
        Q0_CLK1_GTREFCLK_PAD_P_IN       =>      Q0_CLK1_GTREFCLK_PAD_P_IN,
        Q0_CLK1_GTREFCLK_OUT            =>      q0_clk1_refclk_i,
 
        GT0_TXUSRCLK_OUT                =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_OUT               =>      gt0_txusrclk2_i,
        GT0_TXOUTCLK_IN                 =>      gt0_txoutclk_i,
        GT0_TXCLK_LOCK_OUT              =>      gt0_txmmcm_lock_i,
        GT0_TX_MMCM_RESET_IN            =>      gt0_txmmcm_reset_i,
        GT0_RXUSRCLK_OUT                =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_OUT               =>      gt0_rxusrclk2_i,
        GT0_RXOUTCLK_IN                 =>      gt0_rxoutclk_i,
        GT0_RXCLK_LOCK_OUT              =>      gt0_rxmmcm_lock_i,
        GT0_RX_MMCM_RESET_IN            =>      gt0_rxmmcm_reset_i,
 
        GT1_TXUSRCLK_OUT                =>      gt1_txusrclk_i,
        GT1_TXUSRCLK2_OUT               =>      gt1_txusrclk2_i,
        GT1_TXOUTCLK_IN                 =>      gt1_txoutclk_i,
        GT1_TXCLK_LOCK_OUT              =>      gt1_txmmcm_lock_i,
        GT1_TX_MMCM_RESET_IN            =>      gt1_txmmcm_reset_i,
        GT1_RXUSRCLK_OUT                =>      gt1_rxusrclk_i,
        GT1_RXUSRCLK2_OUT               =>      gt1_rxusrclk2_i,
        GT1_RXOUTCLK_IN                 =>      gt1_rxoutclk_i,
        GT1_RXCLK_LOCK_OUT              =>      gt1_rxmmcm_lock_i,
        GT1_RX_MMCM_RESET_IN            =>      gt1_rxmmcm_reset_i,
 
        GT2_TXUSRCLK_OUT                =>      gt2_txusrclk_i,
        GT2_TXUSRCLK2_OUT               =>      gt2_txusrclk2_i,
        GT2_TXOUTCLK_IN                 =>      gt2_txoutclk_i,
        GT2_TXCLK_LOCK_OUT              =>      gt2_txmmcm_lock_i,
        GT2_TX_MMCM_RESET_IN            =>      gt2_txmmcm_reset_i,
        GT2_RXUSRCLK_OUT                =>      gt2_rxusrclk_i,
        GT2_RXUSRCLK2_OUT               =>      gt2_rxusrclk2_i,
        GT2_RXOUTCLK_IN                 =>      gt2_rxoutclk_i,
        GT2_RXCLK_LOCK_OUT              =>      gt2_rxmmcm_lock_i,
        GT2_RX_MMCM_RESET_IN            =>      gt2_rxmmcm_reset_i,
 
        GT3_TXUSRCLK_OUT                =>      gt3_txusrclk_i,
        GT3_TXUSRCLK2_OUT               =>      gt3_txusrclk2_i,
        GT3_TXOUTCLK_IN                 =>      gt3_txoutclk_i,
        GT3_TXCLK_LOCK_OUT              =>      gt3_txmmcm_lock_i,
        GT3_TX_MMCM_RESET_IN            =>      gt3_txmmcm_reset_i,
        GT3_RXUSRCLK_OUT                =>      gt3_rxusrclk_i,
        GT3_RXUSRCLK2_OUT               =>      gt3_rxusrclk2_i,
        GT3_RXOUTCLK_IN                 =>      gt3_rxoutclk_i,
        GT3_RXCLK_LOCK_OUT              =>      gt3_rxmmcm_lock_i,
        GT3_RX_MMCM_RESET_IN            =>      gt3_rxmmcm_reset_i,
        DRPCLK_IN                       =>      DRP_CLK_IN,
        DRPCLK_OUT                      =>      drpclk_in_i

    );

    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    gtx_quad_no_buffer_init_i : gtx_quad_no_buffer_init
    generic map
    (
        EXAMPLE_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION              =>      EXAMPLE_SIMULATION,
        STABLE_CLOCK_PERIOD             =>      STABLE_CLOCK_PERIOD,
        EXAMPLE_USE_CHIPSCOPE           =>      EXAMPLE_USE_CHIPSCOPE
    )
    port map
    (
        SYSCLK_IN                       =>      drpclk_in_i,
        SOFT_RESET_IN                   =>      tied_to_ground_i,
        DONT_RESET_ON_DATA_ERROR_IN     =>      tied_to_ground_i,
        GT0_TX_MMCM_LOCK_IN             =>      gt0_txmmcm_lock_i,
        GT0_TX_MMCM_RESET_OUT           =>      gt0_txmmcm_reset_i,
        GT0_RX_MMCM_LOCK_IN             =>      gt0_rxmmcm_lock_i,
        GT0_RX_MMCM_RESET_OUT           =>      gt0_rxmmcm_reset_i,
        GT0_TX_FSM_RESET_DONE_OUT       =>      gt0_txfsmresetdone_i,
        GT0_RX_FSM_RESET_DONE_OUT       =>      gt0_rxfsmresetdone_i,
        GT0_DATA_VALID_IN               =>      gt0_track_data_i,
        GT1_TX_MMCM_LOCK_IN             =>      gt1_txmmcm_lock_i,
        GT1_TX_MMCM_RESET_OUT           =>      gt1_txmmcm_reset_i,
        GT1_RX_MMCM_LOCK_IN             =>      gt1_rxmmcm_lock_i,
        GT1_RX_MMCM_RESET_OUT           =>      gt1_rxmmcm_reset_i,
        GT1_TX_FSM_RESET_DONE_OUT       =>      gt1_txfsmresetdone_i,
        GT1_RX_FSM_RESET_DONE_OUT       =>      gt1_rxfsmresetdone_i,
        GT1_DATA_VALID_IN               =>      gt1_track_data_i,
        GT2_TX_MMCM_LOCK_IN             =>      gt2_txmmcm_lock_i,
        GT2_TX_MMCM_RESET_OUT           =>      gt2_txmmcm_reset_i,
        GT2_RX_MMCM_LOCK_IN             =>      gt2_rxmmcm_lock_i,
        GT2_RX_MMCM_RESET_OUT           =>      gt2_rxmmcm_reset_i,
        GT2_TX_FSM_RESET_DONE_OUT       =>      gt2_txfsmresetdone_i,
        GT2_RX_FSM_RESET_DONE_OUT       =>      gt2_rxfsmresetdone_i,
        GT2_DATA_VALID_IN               =>      gt2_track_data_i,
        GT3_TX_MMCM_LOCK_IN             =>      gt3_txmmcm_lock_i,
        GT3_TX_MMCM_RESET_OUT           =>      gt3_txmmcm_reset_i,
        GT3_RX_MMCM_LOCK_IN             =>      gt3_rxmmcm_lock_i,
        GT3_RX_MMCM_RESET_OUT           =>      gt3_rxmmcm_reset_i,
        GT3_TX_FSM_RESET_DONE_OUT       =>      gt3_txfsmresetdone_i,
        GT3_RX_FSM_RESET_DONE_OUT       =>      gt3_rxfsmresetdone_i,
        GT3_DATA_VALID_IN               =>      gt3_track_data_i,

  
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X0Y0)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      gt0_drpaddr_i,
        gt0_drpclk_in                   =>      drpclk_in_i,
        gt0_drpdi_in                    =>      gt0_drpdi_i,
        gt0_drpdo_out                   =>      gt0_drpdo_i,
        gt0_drpen_in                    =>      gt0_drpen_i,
        gt0_drprdy_out                  =>      gt0_drprdy_i,
        gt0_drpwe_in                    =>      gt0_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        gt0_loopback_in                 =>      "000",
        ------------------------------ Power-Down Ports ----------------------------
        gt0_rxpd_in                     =>      gt0_rxpd_i,
        gt0_txpd_in                     =>      gt0_txpd_i,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt0_rxcdrlock_out               =>      gt0_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_i,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxdisperr_out               =>      gt0_rxdisperr_i,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_i,
        --------------------------- Receive Ports - RX AFE -------------------------
        gt0_gtxrxp_in                   =>      RXP_IN(0),
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gtxrxn_in                   =>      RXN_IN(0),
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt0_rxphmonitor_out             =>      gt0_rxphmonitor_i,
        gt0_rxphslipmonitor_out         =>      gt0_rxphslipmonitor_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt0_rxmcommaalignen_in          =>      gt0_rxmcommaalignen_i,
        gt0_rxpcommaalignen_in          =>      gt0_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_i,
        gt0_rxpmareset_in               =>      gt0_rxpmareset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt0_rxcharisk_out               =>      gt0_rxcharisk_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt0_txpostcursor_in             =>      gt0_txpostcursor_i,
        gt0_txprecursor_in              =>      gt0_txprecursor_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_i,
        gt0_txuserrdy_in                =>      gt0_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                 =>      gt0_txusrclk_i,
        gt0_txusrclk2_in                =>      gt0_txusrclk2_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt0_txdiffctrl_in               =>      gt0_txdiffctrl_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                   =>      gt0_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gtxtxn_out                  =>      TXN_OUT(0),
        gt0_gtxtxp_out                  =>      TXP_OUT(0),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_i,
        gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_i,
        gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_i,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt0_txcharisk_in                =>      gt0_txcharisk_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt0_txresetdone_i,


  
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X0Y1)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpaddr_in                  =>      gt1_drpaddr_i,
        gt1_drpclk_in                   =>      drpclk_in_i,
        gt1_drpdi_in                    =>      gt1_drpdi_i,
        gt1_drpdo_out                   =>      gt1_drpdo_i,
        gt1_drpen_in                    =>      gt1_drpen_i,
        gt1_drprdy_out                  =>      gt1_drprdy_i,
        gt1_drpwe_in                    =>      gt1_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        gt1_loopback_in                 =>      "000",
        ------------------------------ Power-Down Ports ----------------------------
        gt1_rxpd_in                     =>      gt1_rxpd_i,
        gt1_txpd_in                     =>      gt1_txpd_i,
        --------------------- RX Initialization and Reset Ports --------------------
        gt1_rxuserrdy_in                =>      gt1_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      gt1_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt1_rxcdrlock_out               =>      gt1_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt0_rxusrclk_i,
        gt1_rxusrclk2_in                =>      gt0_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt1_rxdisperr_out               =>      gt1_rxdisperr_i,
        gt1_rxnotintable_out            =>      gt1_rxnotintable_i,
        --------------------------- Receive Ports - RX AFE -------------------------
        gt1_gtxrxp_in                   =>      RXP_IN(1),
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gtxrxn_in                   =>      RXN_IN(1),
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt1_rxphmonitor_out             =>      gt1_rxphmonitor_i,
        gt1_rxphslipmonitor_out         =>      gt1_rxphslipmonitor_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt1_rxmcommaalignen_in          =>      gt1_rxmcommaalignen_i,
        gt1_rxpcommaalignen_in          =>      gt1_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_i,
        gt1_rxpmareset_in               =>      gt1_rxpmareset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt1_rxcharisk_out               =>      gt1_rxcharisk_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt1_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt1_txpostcursor_in             =>      gt1_txpostcursor_i,
        gt1_txprecursor_in              =>      gt1_txprecursor_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_i,
        gt1_txuserrdy_in                =>      gt1_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txusrclk_in                 =>      gt0_txusrclk_i,
        gt1_txusrclk2_in                =>      gt0_txusrclk2_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt1_txdiffctrl_in               =>      gt1_txdiffctrl_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt1_txdata_in                   =>      gt1_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt1_gtxtxn_out                  =>      TXN_OUT(1),
        gt1_gtxtxp_out                  =>      TXP_OUT(1),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclk_out                =>      gt1_txoutclk_i,
        gt1_txoutclkfabric_out          =>      gt1_txoutclkfabric_i,
        gt1_txoutclkpcs_out             =>      gt1_txoutclkpcs_i,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt1_txcharisk_in                =>      gt1_txcharisk_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      gt1_txresetdone_i,


  
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X0Y2)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpaddr_in                  =>      gt2_drpaddr_i,
        gt2_drpclk_in                   =>      drpclk_in_i,
        gt2_drpdi_in                    =>      gt2_drpdi_i,
        gt2_drpdo_out                   =>      gt2_drpdo_i,
        gt2_drpen_in                    =>      gt2_drpen_i,
        gt2_drprdy_out                  =>      gt2_drprdy_i,
        gt2_drpwe_in                    =>      gt2_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        gt2_loopback_in                 =>      "000",
        ------------------------------ Power-Down Ports ----------------------------
        gt2_rxpd_in                     =>      gt2_rxpd_i,
        gt2_txpd_in                     =>      gt2_txpd_i,
        --------------------- RX Initialization and Reset Ports --------------------
        gt2_rxuserrdy_in                =>      gt2_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      gt2_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt2_rxcdrlock_out               =>      gt2_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt0_rxusrclk_i,
        gt2_rxusrclk2_in                =>      gt0_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      gt2_rxdata_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt2_rxdisperr_out               =>      gt2_rxdisperr_i,
        gt2_rxnotintable_out            =>      gt2_rxnotintable_i,
        --------------------------- Receive Ports - RX AFE -------------------------
        gt2_gtxrxp_in                   =>      RXP_IN(2),
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gtxrxn_in                   =>      RXN_IN(2),
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt2_rxphmonitor_out             =>      gt2_rxphmonitor_i,
        gt2_rxphslipmonitor_out         =>      gt2_rxphslipmonitor_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt2_rxmcommaalignen_in          =>      gt2_rxmcommaalignen_i,
        gt2_rxpcommaalignen_in          =>      gt2_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_i,
        gt2_rxpmareset_in               =>      gt2_rxpmareset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt2_rxcharisk_out               =>      gt2_rxcharisk_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt2_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt2_txpostcursor_in             =>      gt2_txpostcursor_i,
        gt2_txprecursor_in              =>      gt2_txprecursor_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_i,
        gt2_txuserrdy_in                =>      gt2_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txusrclk_in                 =>      gt0_txusrclk_i,
        gt2_txusrclk2_in                =>      gt0_txusrclk2_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt2_txdiffctrl_in               =>      gt2_txdiffctrl_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt2_txdata_in                   =>      gt2_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt2_gtxtxn_out                  =>      TXN_OUT(2),
        gt2_gtxtxp_out                  =>      TXP_OUT(2),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclk_out                =>      gt2_txoutclk_i,
        gt2_txoutclkfabric_out          =>      gt2_txoutclkfabric_i,
        gt2_txoutclkpcs_out             =>      gt2_txoutclkpcs_i,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt2_txcharisk_in                =>      gt2_txcharisk_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      gt2_txresetdone_i,


  
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X0Y3)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpaddr_in                  =>      gt3_drpaddr_i,
        gt3_drpclk_in                   =>      drpclk_in_i,
        gt3_drpdi_in                    =>      gt3_drpdi_i,
        gt3_drpdo_out                   =>      gt3_drpdo_i,
        gt3_drpen_in                    =>      gt3_drpen_i,
        gt3_drprdy_out                  =>      gt3_drprdy_i,
        gt3_drpwe_in                    =>      gt3_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        gt3_loopback_in                 =>      "000",
        ------------------------------ Power-Down Ports ----------------------------
        gt3_rxpd_in                     =>      gt3_rxpd_i,
        gt3_txpd_in                     =>      gt3_txpd_i,
        --------------------- RX Initialization and Reset Ports --------------------
        gt3_rxuserrdy_in                =>      gt3_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      gt3_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        gt3_rxcdrlock_out               =>      gt3_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt0_rxusrclk_i,
        gt3_rxusrclk2_in                =>      gt0_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt3_rxdisperr_out               =>      gt3_rxdisperr_i,
        gt3_rxnotintable_out            =>      gt3_rxnotintable_i,
        --------------------------- Receive Ports - RX AFE -------------------------
        gt3_gtxrxp_in                   =>      RXP_IN(3),
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gtxrxn_in                   =>      RXN_IN(3),
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt3_rxphmonitor_out             =>      gt3_rxphmonitor_i,
        gt3_rxphslipmonitor_out         =>      gt3_rxphslipmonitor_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt3_rxmcommaalignen_in          =>      gt3_rxmcommaalignen_i,
        gt3_rxpcommaalignen_in          =>      gt3_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_i,
        gt3_rxpmareset_in               =>      gt3_rxpmareset_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt3_rxcharisk_out               =>      gt3_rxcharisk_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt3_rxresetdone_i,
        ------------------------ TX Configurable Driver Ports ----------------------
        gt3_txpostcursor_in             =>      gt3_txpostcursor_i,
        gt3_txprecursor_in              =>      gt3_txprecursor_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_i,
        gt3_txuserrdy_in                =>      gt3_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txusrclk_in                 =>      gt0_txusrclk_i,
        gt3_txusrclk2_in                =>      gt0_txusrclk2_i,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt3_txdiffctrl_in               =>      gt3_txdiffctrl_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt3_txdata_in                   =>      gt3_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt3_gtxtxn_out                  =>      TXN_OUT(3),
        gt3_gtxtxp_out                  =>      TXP_OUT(3),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclk_out                =>      gt3_txoutclk_i,
        gt3_txoutclkfabric_out          =>      gt3_txoutclkfabric_i,
        gt3_txoutclkpcs_out             =>      gt3_txoutclkpcs_i,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt3_txcharisk_in                =>      gt3_txcharisk_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      gt3_txresetdone_i,




    --____________________________COMMON PORTS________________________________
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        gt0_gtrefclk0_common_in         =>      q0_clk1_refclk_i,
        ------------------------- Common Block - QPLL Ports ------------------------
        gt0_qplllock_out                =>      gt0_qplllock_i,
        gt0_qplllockdetclk_in           =>      drpclk_in_i,
        gt0_qpllpd_in                   =>      gt0_qpllpd_i,
        gt0_qpllreset_in                =>      gt0_qpllreset_i

    );



    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
process(gt0_rxusrclk2_i,gt0_rxresetdone_i)
    begin
        if(gt0_rxresetdone_i = '0') then
            gt0_rxresetdone_r  <= '0'   after DLY;
            gt0_rxresetdone_r2 <= '0'   after DLY;
            gt0_rxresetdone_r3 <= '0'   after DLY;
elsif (gt0_rxusrclk2_i'event and gt0_rxusrclk2_i = '1') then
            gt0_rxresetdone_r  <= gt0_rxresetdone_i   after DLY;
            gt0_rxresetdone_r2 <= gt0_rxresetdone_r   after DLY;
            gt0_rxresetdone_r3  <= gt0_rxresetdone_r2   after DLY;
        end if;
    end process;

process(gt0_txusrclk2_i,gt0_txfsmresetdone_i)
    begin
        if(gt0_txfsmresetdone_i = '0') then
            gt0_txfsmresetdone_r  <= '0'   after DLY;
            gt0_txfsmresetdone_r2 <= '0'   after DLY;
elsif (gt0_txusrclk2_i'event and gt0_txusrclk2_i = '1') then
            gt0_txfsmresetdone_r  <= gt0_txfsmresetdone_i   after DLY;
            gt0_txfsmresetdone_r2 <= gt0_txfsmresetdone_r   after DLY;
        end if;
    end process;
process(gt0_rxusrclk2_i,gt1_rxresetdone_i)
    begin
        if(gt1_rxresetdone_i = '0') then
            gt1_rxresetdone_r  <= '0'   after DLY;
            gt1_rxresetdone_r2 <= '0'   after DLY;
            gt1_rxresetdone_r3 <= '0'   after DLY;
elsif (gt0_rxusrclk2_i'event and gt0_rxusrclk2_i = '1') then
            gt1_rxresetdone_r  <= gt1_rxresetdone_i   after DLY;
            gt1_rxresetdone_r2 <= gt1_rxresetdone_r   after DLY;
            gt1_rxresetdone_r3  <= gt1_rxresetdone_r2   after DLY;
        end if;
    end process;

process(gt0_txusrclk2_i,gt1_txfsmresetdone_i)
    begin
        if(gt1_txfsmresetdone_i = '0') then
            gt1_txfsmresetdone_r  <= '0'   after DLY;
            gt1_txfsmresetdone_r2 <= '0'   after DLY;
elsif (gt0_txusrclk2_i'event and gt0_txusrclk2_i = '1') then
            gt1_txfsmresetdone_r  <= gt1_txfsmresetdone_i   after DLY;
            gt1_txfsmresetdone_r2 <= gt1_txfsmresetdone_r   after DLY;
        end if;
    end process;
process(gt0_rxusrclk2_i,gt2_rxresetdone_i)
    begin
        if(gt2_rxresetdone_i = '0') then
            gt2_rxresetdone_r  <= '0'   after DLY;
            gt2_rxresetdone_r2 <= '0'   after DLY;
            gt2_rxresetdone_r3 <= '0'   after DLY;
elsif (gt0_rxusrclk2_i'event and gt0_rxusrclk2_i = '1') then
            gt2_rxresetdone_r  <= gt2_rxresetdone_i   after DLY;
            gt2_rxresetdone_r2 <= gt2_rxresetdone_r   after DLY;
            gt2_rxresetdone_r3  <= gt2_rxresetdone_r2   after DLY;
        end if;
    end process;

process(gt0_txusrclk2_i,gt2_txfsmresetdone_i)
    begin
        if(gt2_txfsmresetdone_i = '0') then
            gt2_txfsmresetdone_r  <= '0'   after DLY;
            gt2_txfsmresetdone_r2 <= '0'   after DLY;
elsif (gt0_txusrclk2_i'event and gt0_txusrclk2_i = '1') then
            gt2_txfsmresetdone_r  <= gt2_txfsmresetdone_i   after DLY;
            gt2_txfsmresetdone_r2 <= gt2_txfsmresetdone_r   after DLY;
        end if;
    end process;
process(gt0_rxusrclk2_i,gt3_rxresetdone_i)
    begin
        if(gt3_rxresetdone_i = '0') then
            gt3_rxresetdone_r  <= '0'   after DLY;
            gt3_rxresetdone_r2 <= '0'   after DLY;
            gt3_rxresetdone_r3 <= '0'   after DLY;
elsif (gt0_rxusrclk2_i'event and gt0_rxusrclk2_i = '1') then
            gt3_rxresetdone_r  <= gt3_rxresetdone_i   after DLY;
            gt3_rxresetdone_r2 <= gt3_rxresetdone_r   after DLY;
            gt3_rxresetdone_r3  <= gt3_rxresetdone_r2   after DLY;
        end if;
    end process;

process(gt0_txusrclk2_i,gt3_txfsmresetdone_i)
    begin
        if(gt3_txfsmresetdone_i = '0') then
            gt3_txfsmresetdone_r  <= '0'   after DLY;
            gt3_txfsmresetdone_r2 <= '0'   after DLY;
elsif (gt0_txusrclk2_i'event and gt0_txusrclk2_i = '1') then
            gt3_txfsmresetdone_r  <= gt3_txfsmresetdone_i   after DLY;
            gt3_txfsmresetdone_r2 <= gt3_txfsmresetdone_r   after DLY;
        end if;
    end process;

    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    gt0_frame_gen : gtx_quad_no_buffer_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 48)       =>      gt0_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt0_txdata_float16_i,
        TX_DATA_OUT(47 downto 16)       =>      gt0_txdata_i,
 
        TXCTRL_OUT(7 downto 4)          =>      gt0_txcharisk_float_i,
        TXCTRL_OUT(3 downto 0)          =>      gt0_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk2_i,
        SYSTEM_RESET                    =>      gt0_tx_system_reset_c
    );
    
    gt1_frame_gen : gtx_quad_no_buffer_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 48)       =>      gt1_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt1_txdata_float16_i,
        TX_DATA_OUT(47 downto 16)       =>      gt1_txdata_i,
 
        TXCTRL_OUT(7 downto 4)          =>      gt1_txcharisk_float_i,
        TXCTRL_OUT(3 downto 0)          =>      gt1_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk2_i,
        SYSTEM_RESET                    =>      gt1_tx_system_reset_c
    );
    
    gt2_frame_gen : gtx_quad_no_buffer_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 48)       =>      gt2_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt2_txdata_float16_i,
        TX_DATA_OUT(47 downto 16)       =>      gt2_txdata_i,
 
        TXCTRL_OUT(7 downto 4)          =>      gt2_txcharisk_float_i,
        TXCTRL_OUT(3 downto 0)          =>      gt2_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk2_i,
        SYSTEM_RESET                    =>      gt2_tx_system_reset_c
    );
    
    gt3_frame_gen : gtx_quad_no_buffer_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 48)       =>      gt3_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt3_txdata_float16_i,
        TX_DATA_OUT(47 downto 16)       =>      gt3_txdata_i,
 
        TXCTRL_OUT(7 downto 4)          =>      gt3_txcharisk_float_i,
        TXCTRL_OUT(3 downto 0)          =>      gt3_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk2_i,
        SYSTEM_RESET                    =>      gt3_tx_system_reset_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

gt0_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt0_matchn_i;

    -- gt0_frame_check0 is always connected to the lane with the start of char 
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
gt0_inc_in_i                                 <= '0';

    gt0_frame_check : gtx_quad_no_buffer_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      32,
        RXCTRL_WIDTH                    =>      4,
        COMMA_DOUBLE                    =>      x"04bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"060504bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt0_rxdata_i,
        RXCTRL_IN                       =>      gt0_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt0_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt0_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt0_inc_in_i,
        INC_OUT                         =>      gt0_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt0_matchn_i,
        RESET_ON_ERROR_IN               =>      gt0_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt0_rxusrclk2_i,
        SYSTEM_RESET                    =>      gt0_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt0_error_count_i,
        TRACK_DATA_OUT                  =>      gt0_track_data_i
    );

gt1_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt1_matchn_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
gt1_inc_in_i                                 <= gt0_inc_out_i when  (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    gt1_frame_check : gtx_quad_no_buffer_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      32,
        RXCTRL_WIDTH                    =>      4,
        COMMA_DOUBLE                    =>      x"04bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"060504bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt1_rxdata_i,
        RXCTRL_IN                       =>      gt1_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt1_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt1_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt1_inc_in_i,
        INC_OUT                         =>      gt1_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt1_matchn_i,
        RESET_ON_ERROR_IN               =>      gt1_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt0_rxusrclk2_i,
        SYSTEM_RESET                    =>      gt1_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt1_error_count_i,
        TRACK_DATA_OUT                  =>      gt1_track_data_i
    );

gt2_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt2_matchn_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
gt2_inc_in_i                                 <= gt0_inc_out_i when  (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    gt2_frame_check : gtx_quad_no_buffer_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      32,
        RXCTRL_WIDTH                    =>      4,
        COMMA_DOUBLE                    =>      x"04bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"060504bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt2_rxdata_i,
        RXCTRL_IN                       =>      gt2_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt2_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt2_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt2_inc_in_i,
        INC_OUT                         =>      gt2_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt2_matchn_i,
        RESET_ON_ERROR_IN               =>      gt2_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt0_rxusrclk2_i,
        SYSTEM_RESET                    =>      gt2_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt2_error_count_i,
        TRACK_DATA_OUT                  =>      gt2_track_data_i
    );

gt3_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt3_matchn_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
gt3_inc_in_i                                 <= gt0_inc_out_i when  (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    gt3_frame_check : gtx_quad_no_buffer_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      32,
        RXCTRL_WIDTH                    =>      4,
        COMMA_DOUBLE                    =>      x"04bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"060504bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt3_rxdata_i,
        RXCTRL_IN                       =>      gt3_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt3_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt3_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt3_inc_in_i,
        INC_OUT                         =>      gt3_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt3_matchn_i,
        RESET_ON_ERROR_IN               =>      gt3_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt0_rxusrclk2_i,
        SYSTEM_RESET                    =>      gt3_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt3_error_count_i,
        TRACK_DATA_OUT                  =>      gt3_track_data_i
    );




TRACK_DATA_OUT                               <= track_data_out_i;

track_data_out_i                             <= 
                                gt0_track_data_i  and
                                gt1_track_data_i  and
                                gt2_track_data_i  and
                                gt3_track_data_i ;














-------------------------------------------------------------------------------
----------------------------- Debug Signals assignment -----------------------
    gt0_qpllpd_i                                 <= tied_to_ground_i;

------------ optional Ports assignments --------------
gt0_loopback_i                               <= (others => '0');
 
gt0_txdiffctrl_i                             <= (others => '0');
gt0_rxpmareset_i                             <= tied_to_ground_i;
gt0_rxpd_i                                   <= (others => '0');
gt0_txprecursor_i                            <= (others => '0');
gt0_txpostcursor_i                           <= (others => '0');
gt0_txpd_i                                   <= (others => '0');
gt1_loopback_i                               <= (others => '0');
 
gt1_txdiffctrl_i                             <= (others => '0');
gt1_rxpmareset_i                             <= tied_to_ground_i;
gt1_rxpd_i                                   <= (others => '0');
gt1_txprecursor_i                            <= (others => '0');
gt1_txpostcursor_i                           <= (others => '0');
gt1_txpd_i                                   <= (others => '0');
gt2_loopback_i                               <= (others => '0');
 
gt2_txdiffctrl_i                             <= (others => '0');
gt2_rxpmareset_i                             <= tied_to_ground_i;
gt2_rxpd_i                                   <= (others => '0');
gt2_txprecursor_i                            <= (others => '0');
gt2_txpostcursor_i                           <= (others => '0');
gt2_txpd_i                                   <= (others => '0');
gt3_loopback_i                               <= (others => '0');
 
gt3_txdiffctrl_i                             <= (others => '0');
gt3_rxpmareset_i                             <= tied_to_ground_i;
gt3_rxpd_i                                   <= (others => '0');
gt3_txprecursor_i                            <= (others => '0');
gt3_txpostcursor_i                           <= (others => '0');
gt3_txpd_i                                   <= (others => '0');
------------------------------------------------------

    -- assign resets for frame_gen modules
gt0_tx_system_reset_c                        <= not gt0_txfsmresetdone_r2;
gt1_tx_system_reset_c                        <= not gt1_txfsmresetdone_r2;
gt2_tx_system_reset_c                        <= not gt2_txfsmresetdone_r2;
gt3_tx_system_reset_c                        <= not gt3_txfsmresetdone_r2;

    -- assign resets for frame_check modules
gt0_rx_system_reset_c                        <= not gt0_rxresetdone_r3;
gt1_rx_system_reset_c                        <= not gt1_rxresetdone_r3;
gt2_rx_system_reset_c                        <= not gt2_rxresetdone_r3;
gt3_rx_system_reset_c                        <= not gt3_rxresetdone_r3;



end RTL;


