`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MTs+dW5n8qsN7YyJLYWGCcWgD+AnrlpE2UFKli2AoQw4KkGyQKBraU1f20x+SawPQVW+G5DlWKif
JWPlThKA4w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
guMvgNAtq9Ut+YN0I/3BfI+vtSYgU4+vGMAPrVz6r3IUX857KWazizgR/wzf1XwMn6dgl8Hg/wif
3hHdxEH+8k0/6z+6QSKgnaAfaPFnoFYoEtYFVdIQxufP4mIfuVZYWztRJFHPKEtODMhwoEM4wZgH
BwezMe2V+GU8qEh+Eko=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aVYEe2nQzUEKB66PGiEt7bVn5uF3XMZuHAJejzhUbUls6Km4KYttHnegJC5ibGYyyY2wO/dbZ5QG
No5LPds79R/veNIi3cVdguZ42lT41AbjxOFXj99k7e+tL1nDrP/z/K0MXcHsCOAlen1tkN1VxGF6
w7vzK/XxCS2GJlqLDr0uVfuAsZubdo7++lttaRHehY0Llijec1AOl0vvz53Dh6dXeykyHc+RvvJz
Bu0Ktm6+NlSURtWwf3Kq9ZVXd9H+tDYxaDMD9uHjVRgV67fm80WQx1rvgLLHye8UxAZu9usURTwo
CJYlHAe0tIggmUDvmVJsYdI/A9UaGxQn3K7BWw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c+Jc7mg30GoOsKfdrHsqmVtnchPq79zqqREHcqyG7qqc3kcxtNZ3hm8nsOMIXdDv7oY6YFdMjkoY
A6Cu3xlj8R7f+mq8zqZVtjFCnqSbYM5bw3Np1L9dkHv96qy29Ptoi3NJ0iMYfw9XMY8pwOz4bh6y
lJ4wJm07scVUfMv1H94=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rQX0KTjluiuJ8C5MmekfJmaFNHrM4FkUPOKmsRa1CWR2vlrfGQT8cYepWczvHWwTiMcASGB53Aif
tMTJNIRr1dQIYsz1YgY9SCnp3HYGfbDm59RN2kJ5JW4rZ1YADa1ngbvm9aGfYprX+ziMwr4ekThg
UAtD1c+X+qlrPsR1s7ZHDT5JMmeSsYlEaYFq9WVpl7kpU8HSL8a99ZGbhX+YaU+OpRsxP3+BoQ2X
KoQkUhpLW0A+GuTc3U5xsZtBZdHvs9qcoz6zsUjxNAqvgzaLY05c1/eary4B0S3e2pt6BI6ewIbF
SEVb5jBux+G1zuz+kYtf4zyg2aO8rSjyNmbNIw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5664)
`protect data_block
maucsIn9gs8UnRI6PBwXxdHR46caqBfw61uz5teqVuPMi1KD/XvaOqRnAyyXaTYQ/KgpMtoiUOG9
iCH/tYt1SaTuC4RVyh93t/mgGrmE1obJ5bFU5JY9a+GkjRcU5900eid7lGX8jfSfMtcwxiQY0Fxv
VQhkbMxk+UEKt2L93vd6Su5R9TFikdNJz3H1PpPBIZ6tNPtFzruPY+tzYZIFuFjhMGhP2OiEDJZA
xB/yKcGpNg6LD4xm/X3R3gm+ig3MAjUREWAmzLxhs+7meguKXxY0+maF6hcENv4Hen6B9JuJ9DxL
Hxnjh8T66vpRGvzlqQkFG624IGo4oCqWkRT4igddha97OUapgQZY0KlSkLH5OARIlqD8GYlFmwo0
ojBDp+pvdgoMH5NYc2Ut3EUa/2EP0QnJ9ZCHgl7stO0yopUGYPLHzLJYDVQGzy2Lz2gV4j8anQb8
hb+tvfsA9RoHzqlKCX8IX0m2FmlpFzxR4P5ux/SZhlGeZC7FIMz9x1Moo5NT8O3+eDClndeEz8SR
xB/Q4aZfj6sVAmvN7qcpCbEsV6IJb2w3InQu+OPPOIeF3SdVC82xOf5f/DNoUFWq1m8b3xAWWfoy
QHqwBZ0He49i7nB763vCNd+ItJ+bxP4kJ3ntYRfdc0502eVKxGE+cB/GMY6QFUHXh3Ikhn5nSCFf
0Ns7/A4ROocGy8kLhM6fgpJRSKYP11Quic7hJXpkdc1eN5OOTEqaoKudUoqDmyKl+e4g8UO2xn0P
qLFj6FtyJgydA9fmvctMUCuRZ0Q+VZ0VdzfMWayDSw56oA0FdoV4a5Hkkd3BNNqL6hsy5Om9R+DW
Hf0YGtzksfDzXdfRpIbaAlD8oyO5FXnrLG/2F7hLU1z5fQUn4x78fXrhdtNz0wbD0D/JvX5t3RxU
1cSGvAl2gjuNWbAPRYP8SgYGp8UmfH0IFrQpHDNZnW2I+XAK4xJHeAO6rqEYrRxlJ3k7gJpAlqgU
KzjtXXEP6w1J+XGhQUZkrBWoNELvALteB3/V5SoA87oWZ1CrmFnMNWsYV557RlJAK1FhhEhThi+e
Tf3tsubEdKoxkQNhkkNlb/E5/OFEAVQmOdRmE6jcCOz5wfdu57nouk/TeflBE5rU49AXZFeN0MRG
bFV5hm897JQy7xFHtLAp7Kj2By5YkE8NN1myOPeIAoix4qrpTSxr6V8sWhyfdEPakeB/n/crXhwq
POvVakvuJFXaIZouJAJnSjGqzjhpc9Or+NyQA7MqhBUgPyvE5VxDDmArCe/wDLC0ja2FDHjTv/xT
Ofnhv8vWnNrKX76FNuJCGRnFgiGnsboHUujQRKcDH/5EkqVBeuUSFz5QjdLlZdt19PE+54DEBmMr
8OhVPwOpUk5DxD4nHOMxoHzDuEWVRfHq6tnVxdHRrav29WP8XFRjtfHhLXR2vexPqkaU+9XeJzKl
1Wfm4Gbl0TrenegrLJRzJgTV+nrb6w26YD3qFzc8/GE0dRJytVkdM4UFCRDOIcbKwRisFTamhGIh
iK0e4fwJbmsEaw9rkTB4TxV9MzfN6/aPumad7Iuin6GzcMRVWxirFQtMy1uqXNiLF3YRTWoxFxd8
y7VIbPNhyNlA6kX1C0/U/u0lHGSS7zU3B1F9RK8uTGRte51msSAqYSkmHzM3a2GBhjlIT/ipQkLN
bwlWlheJj3dUO2OWrAF17KKuQbGnryEOjmOqlZ2vCeMU7mHSoBeQNAWsQGPS1ZNoxwTMyDnwLchO
BSN4tS3tkCF2N91d7ooxAqoNAl704MQhXC8f/2BRK1dD2zUL7JcC/NRZ7oKpi/uDTi2Pt6MwC0wk
J5e1FU8k7xnRe1sVf4oaYQwN+KfvkbvZ74cY7S9PA4v8HoplhewgCsFuFlyABTpCisQ5/ZIqdMVa
HBKHup569b6LCxpEwG5py/Uy7fsyIM0v0PULh1BtzsEsQfXf7CD4apuRUr6+F1bip2uOm4zveP70
nQRY0cQqvaLW3aQkJZy5V2F5ZUccI75zTasaaKEcfeFwylBGOz+lkEy58pcixWgpvTtPRDtET/Zr
g6lKtG3SBh3Ug27DxA18hl/ZFuT0FHfVN7544MecfXPJ4oFbFxzLru1xsSlRgFFdF//OKG0S3L67
ypxxgUnZCceU0n9nBhkr/5acuuDXCy+lMZ0Ng0eHfI3ChVvc1ZFdmBhf+dZnDUZm5btKkbaxPzGM
Vr1DwSKTkwzW2AcPHLPo3adURFWR46IDGZnLd1fg5zzswHsqC8BgNuW4AfSOfAZp+t9Huk9k/LJu
DeZOaeJkaTzBjQwrzk2vZ4Y6P6X1uj2H8158jx4Cg0Ahct7ZnLc1JeX0w5qHnckd6MgA+61jMkc7
8JgNWOhunqe1E3JPDCoTjNOStzbRYx36pDXRI2a9e3RwnmZF8C60FPdEqz0zEsvdnm3HhXO8PuYB
kToVB3gGtfsqEh8mwtq9CRyYHRwQcofhZ7gNZVAF1kxttKbHmoYA/HbY2Z1EqaThnkOpes4Sw0AY
C/lhlVxUEfLcoAOwrUBMfTOflDSAlkW/dmjvFJwMyp3kSk3H3Ac3NMutIZPoPLEDTh7rRVaOeAcv
8FEod8WVg4t/r9FstGpAtyUWv8RvQbl/c9o2GZIsO8FM2pNFg66sfbdD2rAZYPnyVPg+tuY89uKm
Gf+4FjCS0HDbh8ywM6yxJRsD1JDIqoNS5jyZp4Kz0LAsFnAf+0KCPmTdn+hUTmBdMRXKKtMSFq7+
9ykOQolgVyXKE8plujYZ1Icdqi+LW1jJOy+STR0MGvr5pDd7QQTQXo837hlVpA+3ZJEDmVuO1+Lu
j0HRDd2laEswkJnvpDnnTi6hFtdnMUW5GgY34zgyETRYyMNLiKi1Gkk6pq5m6zyYrFZAWve5SBO2
fLRf2itBmJiOPNikcDwRYWR5R6XoLOabhKiwbPEUFdgTNxTTURvqg441mYdYwMgXfEWha9Iy1ggf
yONZ99qXfNAhzzXGehudrbQrwcsxKv3SQEl1BSZuwkNRh3k1azUcZYFUoIJwRvjiMakJy50N32du
iRGwI4Lt4NiFdwsXBGjUsR0XauvSt4e9DX34HdcjhVCwWV4EjMVZ/tDft8DZnuzwVGqNrjEHMeSL
tGa2fwUh76PvCi+BUd6Kz4VHyQoxKxeY8CLjRd3VVhzcJwnnujyqAKd4yINvtv8u6+BjEF06og0o
S/SiBX5c9ASwJUI+uyBGQY35FhJJ/6AtHeRMNXUI2gbdUFqS3frIjtYXV7l/jcz0NkVvhKQ9jA99
nGDYmvQYi2vGU5crC+2yCAOZLSCvwpm3ED+kWBsJCTLTsIkEkPpKkpIRbzT4G/jE+Z2NZrMu77+l
44StikvwCg022HmAWseelbyoNInsfAMRACM0r76W+JEQdiNJdqs7to/q9UVCgLZQl41/6SOFpAzq
8xIlK/iw15tuRiGqm6a1rGAHjhL2cXVcvDmomVESxsruNV4ae6eN3H1T0uk323P7Y+Xlzqfoaxdv
oVOPE+iCT/+5CsR1z/f2qt++YEe9ekI+qabaLaSfAdGbDCll7tDe9rUEI5IAJk0b70nzX7eO++fG
ezWPFzFP98TflHYxa6AjA2HF3dKuWLWjh2rSK2c3KGB4UVs0/KhWGPit6mdAujfkdiooWpWATGN5
99cKY1VYNtDtLDsYG4GQ466bwUczXb+ut1jp98+1TXKo3F6Epb6rWKHqCKlmHYfvRa0+zfamH2S5
e3HuBhNEA+WpAPbNTV9pAeoIFKR1CE5Yj6xDWpXi2RGnD0M6QKBqkLo2f1aqDLuyWNyGvC8l8u3M
Z5E/6dvrFSCvoaqTFGPLhKoAdoMzt7tRIqWEj536/3ORJky/yDV4YA9N0R3PPLnDBoFUj70Q6O0t
mzgwev/Z9ONN8dQu7K6jSSZxPAsevyZXgAbYJS9dbPwEj0mcm4OQCbsNscAljJ3AkBF8hdMr/y4z
dKxtAUqSo62HPEr+RbLEf6fO72kI58bVqEIJaHYUJBONArTiNMEIONt+ptvWta8MqRIHftLY4Tyu
wxFnIm8RPYJEpsT89BChvwXRtYDth2QcghAd1ENXAghSzy+k7KJWLeMMJg1d45Xhs+DQY3YMzhwa
kGYDm2AahLrTLwmttE9y+SiUr5NP3C4oZxYKPjA6LQZ4sL6Duq2jjQiYH4KlcI8vs33x3p1xF/8x
+cytgaTwXPhCx0xRcXteGB6Z2obMQtk7koTW77LX7t6lPBxJdlL+CCnTiMkMUeOxfOAQjKRTHlk4
t64LlhtDk+tAd8tFb5w3tIQqluvoR/SNe8mqnWz/ZQCgwKVDAieaPCG85P/z5kgWpBE16qumcA01
VYIL/JftDkSOW4BZfNSKxQYvxEoTehjl4pR1ilMgZNiStMh6sLgX+nUag3w83c8b44PdLHbzCYVB
AUS3gVY3W8t0t09BPF5pPW4FDUpU6X106pKwJVM8E8T8RZGHehb8/iUqlAQhKPLoBEELu1L0KbEu
25WeG/OW0dzYHpFP7DrMpYsRSw0/KiHn4mAxW6ozU6gy03rE7depNMHXqDMb0FghDMRUP1OY5K3/
pAHlQn30rCFlzInxeBEfQlyfPe50k8hODdVwtbgilbD0FQE5MBpcikeQdLwxlVHXtkhqQBgwoHsE
ZZxr0EDYzL21+5Dfbv5VthEM5X/TPYiGAzYC36lD0NCPR51yXyBe7BezQaBludHv9L57BD6kfPAt
tVVgAFUjBJAqFbGTs5k/oQTQKdxzx+pD24mWoLU+r6VEXrqn0tDUp9l/zqWUQ66jdTId8v+VcLiq
nxlCZq1eQ4e/nnaTZY2XQC8OgUMGP3XXdm30MqwhjW8pTaQWDzTwR68yDrbUBz6NDlwBrmi1AqSx
har7tz2AmOKyrV3U38P+Ab3NMuQSkwcSaMS9ncqsCAEaA9rxFzoDyby4cPRhIHM+6BlJeHBFr28e
JpAd02xQ/8lMioZ+OYbS+ZAsb2DTeZSoJYMXJeIUIy40jKGaja7LINk8lEhh6TNMFCwjFRId4acJ
5N+hgU4HDPMQG/VsgOpwzMg91bfoYbCJLI7lurFhsSXdJzqRDdE9BkqCMp5L3Pf/F9Jz2/OC7cPL
0K5avg5s9w9F8eOcNiHmXKO9VWKqEiqhenz4+RjMP3YK5k050KXMaFIdJMGcS3QiUP115jxglxnB
R+n7MahObi88XelhKcumiZxW5Kjfm+aHb7CFs8fs2e+8U6iU95IfmPtAu2TB6Oh0cOPSfNkXSwbM
yvA3iWnRZKEkADD6+RSLUEQuxiDE3V8ANAqCrZkNo2JfEWfj02UbwaeF3jeTE2viXxZKxAXtpWyz
vOfBPXOFBGkDuSzgEhOm/jNKyCziNlCo4s/+X/LpDdBXcLQVMAyTaaj1xRkobSa7P8hiI9v4H768
z31aKjwvUv6t0VCcR+BQZ2Pa6EnKR8sl99uuqjemwc+RUad7LR+2F/NYG6D9iLBPN9qc3pSOjzB8
II9AYw5O769AV4yVwSFQMo9Q8UPZFhGLs12jZcVC5QOhJN5Qox327RFMezqbo5WSwvF5JayCaY5u
g9EwcnMRxXIpUMhXmWUqKbHSoeks7FwZD6owYlBa5D8XOM/5/hth6tHKPs49I7dtZV9xbNIaLBKe
sM2KYp4AI1Gg+wuGPFL3g9IQa3XfDnVTpftOw7CC8BmI2TbWDFk37SeAgxBYXLRoG+WeNa0kvfuF
H3kSptgLTyC65eXk/u5t269R9fQLPy31+v2PDnpA0gj49N9DcyPw7Hmhujnt7nWFUNZEoQ0XqhPh
ZWANsSItE/jBw0rbJnORTF28TXmmBHaoxJ9wLsrvCxjAVBpsa8u1hKRtdNQuwl4JuQWhBvMAWAtD
vxIZCkKUO7OjCd8CKk3kYV/w6ofeCViJ259Kyarh1LR2Xr59XDOOGdhK+ceyROBdNXPi3cHOiSLL
1xBLjEe08ImjaJ1otggNZ/lBI2vXlkBEwbNRTyyXLAA+YBy3ocn127ISn502kBfXXt0wHl4jyi1V
iio5UF+vZD8vZrAhjuDPxizeSvDH/EGQ/f3BtkeHXJ52jPdiYpCipjkg8IFc/LdYF3jNQhXb1Jwv
rFQehlCvqRzNTD21enWb6166ldGsEFgh5f8A2Ru9GVyPt3GkBvQXIvj9g/rEF1txG4bOup7BTG7b
UYVrFg9jQFEGj9vLVbYnrzLvJ2z8/YTrRusoC1qPJdDoN3IhPSj/LsOgMXU+gvviXPbB4rQBVRiO
7g8pGzqqjrQr4nPbaNEe0GRv1lDOmNmDY5yirL0B27DW3b20io3U6+mba1TNSMpeDg9JF+g539AX
R/7mrhGG2qxH5LzGthXghUU48Tr0uhOa/H4H7y4stJq4weFOv9RLsrv1eHDW7pnj4pnI/J84ZvYz
e2+neYqYIcJ6EuD9LRNEiGgbxQnrEcD/OA7JPlDVsMaxdN6PoB5NSh3qZ0dxN2T7amTkGWRryISf
+l8Wb9GDEzdtJwxw+KWMa4NXhC7LE/8eJizuaGN7xedKUooN7vY39Fcvi4NUTkzyFwtFLPDm44Ge
GsyGoNVRWrkRujMp8ZTqmMARNcFEe+PJMgD/eWwYTUdfF/JU37VTaEX88RaQCavR0WESX8c0B5H2
IgCZ+QuxgVEPQgFPbAZzPwhKdfnGCWmSOwDMZjUyCJsi9/zoLjoZb07rtsGwWjEI2aF4KR09GoXc
8joL4qrsmTdZdJTOlYfUtOdHInVxOxFeOqcQA4bGl7ZNNpmfESaVI8RMgZAvCCHazAnVrRUiT5Z0
6Fq0/kGqIzT8sLqBBX1+kdDMbM90p1dqkGghfIg2mDmXL42V1aAfUmM5SmX8EtlHVPCBhn2xa0Ow
EKvZNerOeUmIlr7AqxYWCGeMk5kMKkbos1kQQyLXYfwX2H9ibAF5AxEUu4EzvP84XFKb0V5m2qxw
xeyU2pc9L0gWG5Z/xUeeyi+gUdyD7MMeLF+JI2FxIEHy/5jkI7dqWF1wRRWJN6z/pwOPRAn3GLHS
J4o7JfMiAKqhEWLCdJvhbqZ1WMtOiK33bIp0Znf/lhtz3K29A7z/yvhoB/DK7pUZ9dTi4JQejaqx
ugrYSoWakkiu9jOgCpvEV9wM5tc+E9iDZ9rCXjw86fa5LeBrNiCsAucJkHdKjgwrS1XBYOwawuU0
4y59koT+zGr8ueY3EjgOnVCVK0WL/P82u7QGDICBIP/ZRIQceOSks/EWV0bNxS08k1UX+oJeXcu5
ZVthu3GliAdiF6zxb70euFPtp+TIXPYYwicgOisci5SCy1P81hk5YrX+oFyBeemv0Quam4Poe8og
20I4e8UrQGyP//J+gObAyLP9W8wZpLV0/LP6wR8f4s1NpPtJOWPVFp50bPUwnU2jeL/lMP6PbFCh
02c8WYBpyEtSIBjIKWrkl/+wEFCWzCxwjZkBPhTqte7n7mC7mplkEnLiU9In1q7gb6qrTl5QxgZY
7PQHnnH60QyCgSbEHp6tITOdX2a/OA/bo1z5sLRzUTUe8CSBRvsDvS4rku6g6vqr7UUijyzY8UMT
bZ57yeAuXXOgDb/gc4qko72irpk+
`protect end_protected
