library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.L1TopoDataTypes.all;

Package L1TopoFunctions is
	function ld(m : positive) return natural;
	function sqrt(d : UNSIGNED) return UNSIGNED;
	function reg_ctrl(ctrl_reg_flags : std_logic_vector) return integer;
	function find_msb_1(input : std_logic_vector) return integer;
	function calc_crc(data : std_logic_vector(115 downto 0)) return std_logic_vector;
--	function Jet_TOB_to_std_logic_vector(arg : JetTOB) return std_logic_vector;
--	function std_logic_vector_to_Jet_TOB(arg : std_logic_vector(27 downto 0)) return JetTOB;
	function std_logic_vector_to_TOB(arg : std_logic_vector(22 downto 0); phi_bit4 : std_logic; phi_bit5 : std_logic) return ClusterTOB;
	function std_logic_vector_to_TOB(arg : std_logic_vector(21 downto 0)) return GenericTOB;
	function std_logic_vector_to_TOB(arg : std_logic_vector(27 downto 0); phi_bit1 : std_logic) return JetTOB;
	function std_logic_vector_to_TOB(arg : std_logic_vector(7 downto 0)) return MuonTOB;
--	function TOB_to_std_logic_vector(arg : ClusterTOB) return std_logic_vector;
--	function TOB_to_std_logic_vector(arg : JetTOB) return std_logic_vector;
--	function TOB_to_std_logic_vector(arg : GenericTOB) return std_logic_vector;
--	function TOB_to_std_logic_vector(arg : MuonTOB) return std_logic_vector;
	function to_GenericTOB(arg : ClusterTOB) return GenericTOB;
	function to_GenericTOB(jet : JetTOB; jet_size : integer) return GenericTOB;
	function to_GenericTOB(arg : MuonTOB) return GenericTOB;
	function is_in_eta_range(eta_bin : std_logic_vector;
		                      min_bin : std_logic_vector;
		                      max_bin : std_logic_vector) return boolean;
end package L1TopoFunctions;

Package body L1TopoFunctions is

	-- log_2 function
	function ld(m : positive) return natural is
	begin
		for n in 0 to integer'high loop
			if (2 ** n >= m) then
				return n;
			end if;
		end loop;
	end function ld;

	--sqrt function
	function sqrt(d : UNSIGNED) return UNSIGNED is
		variable a              : unsigned(31 downto 0) := d; --original input.
		variable q              : unsigned(15 downto 0) := (others => '0'); --result.
		variable left, right, r : unsigned(17 downto 0) := (others => '0'); --input to adder/sub.r-remainder.
	begin
		for i in 0 to 15 loop
			right(0)           := '1';
			right(1)           := r(17);
			right(17 downto 2) := q;
			left(1 downto 0)   := a(31 downto 30);
			left(17 downto 2)  := r(15 downto 0);
			a(31 downto 2)     := a(29 downto 0); --shifting by 2 bit.
			if (r(17) = '1') then
				r := left + right;
			else
				r := left - right;
			end if;
			q(15 downto 1) := q(14 downto 0);
			q(0)           := not r(17);
		end loop;
		return q;
	end sqrt;
	
	-- find number of "1" (from right side) in ctrl_flags
	-- TODO: Check if it works correctly!
	function reg_ctrl(ctrl_reg_flags : std_logic_vector) return integer is
		variable ctrl_flags : std_logic_vector(ctrl_reg_flags'length - 1 downto 0);
		variable result     : integer;
	begin
		ctrl_flags := ctrl_reg_flags;
		result     := -1;
		for i in 0 to ctrl_reg_flags'length - 1 loop
			if ctrl_flags(i) = '0' then
				result := i;
				return result;
			end if;
		end loop;
		return -1;
	end;
	
	-- find most significant bit set to "1"
	function find_msb_1(input : std_logic_vector) return integer is
		variable temp       : std_logic_vector(input'length - 1 downto 0);
		variable result     : integer;
	begin
		temp   := input;
		result := 0;
		for i in input'length - 1 downto 0 loop
			if temp(i) = '1' then
				result := i;
				return result;
			end if;
		end loop;
		return 0;
	end;

	-- calculate crc data
	function calc_crc(data : std_logic_vector(115 downto 0)) return std_logic_vector is
		variable d       : std_logic_vector(115 downto 0);
		variable new_crc : std_logic_vector(11 downto 0);
	begin
		d := data;

		new_crc(0) := d(0) xor d(8) xor d(9) xor d(10) xor d(11) xor d(12) xor d(16) xor d(18) xor d(20) xor d(22) xor d(25) xor d(28) xor d(30) xor d(35) xor d(41) xor d(42) xor d(43) xor d(44) xor d(45) xor d(46) xor d(47) xor d(49) xor d(51) xor d(53)
			xor d(54) xor d(55) xor d(58) xor d(59) xor d(61) xor d(62) xor d(64) xor d(65) xor d(66) xor d(67) xor d(69) xor d(71) xor d(72) xor d(78) xor d(79) xor d(80) xor d(81) xor d(84) xor d(86) xor d(88) xor d(91) xor d(92) xor d(96) xor d(100) xor d(
				105) xor d(106) xor d(107) xor d(109) xor d(110) xor d(111) xor d(112) xor d(113) xor d(115);
		new_crc(1) := d(0) xor d(1) xor d(8) xor d(13) xor d(16) xor d(17) xor d(18) xor d(19) xor d(20) xor d(21) xor d(22) xor d(23) xor d(25) xor d(26) xor d(28) xor d(29) xor d(30) xor d(31) xor d(35) xor d(36) xor d(41) xor d(48) xor d(49) xor d(50)
			xor d(51) xor d(52) xor d(53) xor d(56) xor d(58) xor d(60) xor d(61) xor d(63) xor d(64) xor d(68) xor d(69) xor d(70) xor d(71) xor d(73) xor d(78) xor d(82) xor d(84) xor d(85) xor d(86) xor d(87) xor d(88) xor d(89) xor d(91) xor d(93) xor d(
				96) xor d(97) xor d(100) xor d(101) xor d(105) xor d(108) xor d(109) xor d(114) xor d(115);
		new_crc(2) := d(0) xor d(1) xor d(2) xor d(8) xor d(10) xor d(11) xor d(12) xor d(14) xor d(16) xor d(17) xor d(19) xor d(21) xor d(23) xor d(24) xor d(25) xor d(26) xor d(27) xor d(28) xor d(29) xor d(31) xor d(32) xor d(35) xor d(36) xor d(37)
			xor d(41) xor d(43) xor d(44) xor d(45) xor d(46) xor d(47) xor d(50) xor d(52) xor d(55) xor d(57) xor d(58) xor d(66) xor d(67) xor d(70) xor d(74) xor d(78) xor d(80) xor d(81) xor d(83) xor d(84) xor d(85) xor d(87) xor d(89) xor d(90) xor d(
				91) xor d(94) xor d(96) xor d(97) xor d(98) xor d(100) xor d(101) xor d(102) xor d(105) xor d(107) xor d(111) xor d(112) xor d(113);
		new_crc(3) := d(0) xor d(1) xor d(2) xor d(3) xor d(8) xor d(10) xor d(13) xor d(15) xor d(16) xor d(17) xor d(24) xor d(26) xor d(27) xor d(29) xor d(32) xor d(33) xor d(35) xor d(36) xor d(37) xor d(38) xor d(41) xor d(43) xor d(48) xor d(49)
			xor d(54) xor d(55) xor d(56) xor d(61) xor d(62) xor d(64) xor d(65) xor d(66) xor d(68) xor d(69) xor d(72) xor d(75) xor d(78) xor d(80) xor d(82) xor d(85) xor d(90) xor d(95) xor d(96) xor d(97) xor d(98) xor d(99) xor d(100) xor d(101) xor d(
				102) xor d(103) xor d(105) xor d(107) xor d(108) xor d(109) xor d(110) xor d(111) xor d(114) xor d(115);
		new_crc(4) := d(0) xor d(1) xor d(2) xor d(3) xor d(4) xor d(8) xor d(10) xor d(12) xor d(14) xor d(17) xor d(20) xor d(22) xor d(27) xor d(33) xor d(34) xor d(35) xor d(36) xor d(37) xor d(38) xor d(39) xor d(41) xor d(43) xor d(45) xor d(46) xor
			d(47) xor d(50) xor d(51) xor d(53) xor d(54) xor d(56) xor d(57) xor d(58) xor d(59) xor d(61) xor d(63) xor d(64) xor d(70) xor d(71) xor d(72) xor d(73) xor d(76) xor d(78) xor d(80) xor d(83) xor d(84) xor d(88) xor d(92) xor d(97) xor d(98)
			xor d(99) xor d(101) xor d(102) xor d(103) xor d(104) xor d(105) xor d(107) xor d(108) xor d(113);
		new_crc(5) := d(1) xor d(2) xor d(3) xor d(4) xor d(5) xor d(9) xor d(11) xor d(13) xor d(15) xor d(18) xor d(21) xor d(23) xor d(28) xor d(34) xor d(35) xor d(36) xor d(37) xor d(38) xor d(39) xor d(40) xor d(42) xor d(44) xor d(46) xor d(47) xor
			d(48) xor d(51) xor d(52) xor d(54) xor d(55) xor d(57) xor d(58) xor d(59) xor d(60) xor d(62) xor d(64) xor d(65) xor d(71) xor d(72) xor d(73) xor d(74) xor d(77) xor d(79) xor d(81) xor d(84) xor d(85) xor d(89) xor d(93) xor d(98) xor d(99)
			xor d(100) xor d(102) xor d(103) xor d(104) xor d(105) xor d(106) xor d(108) xor d(109) xor d(114);
		new_crc(6) := d(2) xor d(3) xor d(4) xor d(5) xor d(6) xor d(10) xor d(12) xor d(14) xor d(16) xor d(19) xor d(22) xor d(24) xor d(29) xor d(35) xor d(36) xor d(37) xor d(38) xor d(39) xor d(40) xor d(41) xor d(43) xor d(45) xor d(47) xor d(48)
			xor d(49) xor d(52) xor d(53) xor d(55) xor d(56) xor d(58) xor d(59) xor d(60) xor d(61) xor d(63) xor d(65) xor d(66) xor d(72) xor d(73) xor d(74) xor d(75) xor d(78) xor d(80) xor d(82) xor d(85) xor d(86) xor d(90) xor d(94) xor d(99) xor d(
				100) xor d(101) xor d(103) xor d(104) xor d(105) xor d(106) xor d(107) xor d(109) xor d(110) xor d(115);
		new_crc(7) := d(3) xor d(4) xor d(5) xor d(6) xor d(7) xor d(11) xor d(13) xor d(15) xor d(17) xor d(20) xor d(23) xor d(25) xor d(30) xor d(36) xor d(37) xor d(38) xor d(39) xor d(40) xor d(41) xor d(42) xor d(44) xor d(46) xor d(48) xor d(49)
			xor d(50) xor d(53) xor d(54) xor d(56) xor d(57) xor d(59) xor d(60) xor d(61) xor d(62) xor d(64) xor d(66) xor d(67) xor d(73) xor d(74) xor d(75) xor d(76) xor d(79) xor d(81) xor d(83) xor d(86) xor d(87) xor d(91) xor d(95) xor d(100) xor d(
				101) xor d(102) xor d(104) xor d(105) xor d(106) xor d(107) xor d(108) xor d(110) xor d(111);
		new_crc(8) := d(4) xor d(5) xor d(6) xor d(7) xor d(8) xor d(12) xor d(14) xor d(16) xor d(18) xor d(21) xor d(24) xor d(26) xor d(31) xor d(37) xor d(38) xor d(39) xor d(40) xor d(41) xor d(42) xor d(43) xor d(45) xor d(47) xor d(49) xor d(50)
			xor d(51) xor d(54) xor d(55) xor d(57) xor d(58) xor d(60) xor d(61) xor d(62) xor d(63) xor d(65) xor d(67) xor d(68) xor d(74) xor d(75) xor d(76) xor d(77) xor d(80) xor d(82) xor d(84) xor d(87) xor d(88) xor d(92) xor d(96) xor d(101) xor d(
				102) xor d(103) xor d(105) xor d(106) xor d(107) xor d(108) xor d(109) xor d(111) xor d(112);
		new_crc(9) := d(5) xor d(6) xor d(7) xor d(8) xor d(9) xor d(13) xor d(15) xor d(17) xor d(19) xor d(22) xor d(25) xor d(27) xor d(32) xor d(38) xor d(39) xor d(40) xor d(41) xor d(42) xor d(43) xor d(44) xor d(46) xor d(48) xor d(50) xor d(51)
			xor d(52) xor d(55) xor d(56) xor d(58) xor d(59) xor d(61) xor d(62) xor d(63) xor d(64) xor d(66) xor d(68) xor d(69) xor d(75) xor d(76) xor d(77) xor d(78) xor d(81) xor d(83) xor d(85) xor d(88) xor d(89) xor d(93) xor d(97) xor d(102) xor d(
				103) xor d(104) xor d(106) xor d(107) xor d(108) xor d(109) xor d(110) xor d(112) xor d(113);
		new_crc(10) := d(6) xor d(7) xor d(8) xor d(9) xor d(10) xor d(14) xor d(16) xor d(18) xor d(20) xor d(23) xor d(26) xor d(28) xor d(33) xor d(39) xor d(40) xor d(41) xor d(42) xor d(43) xor d(44) xor d(45) xor d(47) xor d(49) xor d(51) xor d(52)
			xor d(53) xor d(56) xor d(57) xor d(59) xor d(60) xor d(62) xor d(63) xor d(64) xor d(65) xor d(67) xor d(69) xor d(70) xor d(76) xor d(77) xor d(78) xor d(79) xor d(82) xor d(84) xor d(86) xor d(89) xor d(90) xor d(94) xor d(98) xor d(103) xor d(
				104) xor d(105) xor d(107) xor d(108) xor d(109) xor d(110) xor d(111) xor d(113) xor d(114);
		new_crc(11) := d(7) xor d(8) xor d(9) xor d(10) xor d(11) xor d(15) xor d(17) xor d(19) xor d(21) xor d(24) xor d(27) xor d(29) xor d(34) xor d(40) xor d(41) xor d(42) xor d(43) xor d(44) xor d(45) xor d(46) xor d(48) xor d(50) xor d(52) xor d(53)
			xor d(54) xor d(57) xor d(58) xor d(60) xor d(61) xor d(63) xor d(64) xor d(65) xor d(66) xor d(68) xor d(70) xor d(71) xor d(77) xor d(78) xor d(79) xor d(80) xor d(83) xor d(85) xor d(87) xor d(90) xor d(91) xor d(95) xor d(99) xor d(104) xor d(
				105) xor d(106) xor d(108) xor d(109) xor d(110) xor d(111) xor d(112) xor d(114) xor d(115);
		return new_crc;
	end calc_crc;

	--------------------------------------------------------
	-- Functions to convert TOBs from/to std_logic_vector --
	--------------------------------------------------------
	
--	function Jet_TOB_to_std_logic_vector(arg : JetTOB) return std_logic_vector is
--		variable result : std_logic_vector(28 downto 0);
--	begin
--		result(18 downto 10) := arg.Et1;
--		result(9 downto 0)   := arg.Et2;
--		result(23 downto 19) := arg.Eta;
--		result(28 downto 24) := arg.Phi;
--		return result;
--	end function Jet_TOB_to_std_logic_vector;

--	function std_logic_vector_to_Jet_TOB(arg : std_logic_vector(28 downto 0)) return JetTOB is
--		variable result : JetTOB;
--	begin
--		result.Et1 := arg(18 downto 10);
--		result.Et2 := arg(9 downto 0);
--		result.Eta := arg(23 downto 19);
--		result.Phi := arg(28 downto 24);
--		return result;
--	end function std_logic_vector_to_Jet_TOB;

	function std_logic_vector_to_TOB(arg : std_logic_vector(22 downto 0); phi_bit4 : std_logic; phi_bit5 : std_logic) return ClusterTOB is
		variable result : ClusterTOB;
	begin
		result.Et              := arg(7 downto 0);
		result.Isol            := arg(12 downto 8);
		result.Eta             := arg(18 downto 13);
		result.Phi(3 downto 0) := arg(22 downto 19);
		result.Phi(4)          := phi_bit4; --!
		result.Phi(5)          := phi_bit5; --!
		return result;
	end function std_logic_vector_to_TOB;

	function std_logic_vector_to_TOB(arg : std_logic_vector(21 downto 0)) return GenericTOB is
		variable result : GenericTOB;
	begin
		result.Et  := arg(9 downto 0);
		result.eta := arg(15 downto 10);
		result.phi := arg(21 downto 16);
		return result;
	end function std_logic_vector_to_TOB;

	function std_logic_vector_to_TOB(arg : std_logic_vector(27 downto 0); phi_bit1 : std_logic) return JetTOB is
		variable result : JetTOB;
	begin
		result.Et1 := arg(18 downto 10);
		result.Et2 := arg(9 downto 0);
		result.Eta := arg(23 downto 19);
		result.Phi(0)          := arg(24);
		result.Phi(1)          := phi_bit1; --!
		result.Phi(4 downto 2) := arg(27 downto 25);
		return result;
	end function std_logic_vector_to_TOB;

	function std_logic_vector_to_TOB(arg : std_logic_vector(7 downto 0)) return MuonTOB is
		variable result : MuonTOB;
	begin
		result.Eta := arg(7 downto 5);
		result.Phi := arg(4 downto 2);
		result.Pt  := arg(1 downto 0);
		return result; -- TODO: Check if this is correct!
	end function std_logic_vector_to_TOB;

--	function TOB_to_std_logic_vector(arg : ClusterTOB) return std_logic_vector is
--		variable result : std_logic_vector(24 downto 0);
--	begin
--		result(7 downto 0)   := arg.Et;
--		result(12 downto 8)  := arg.Isol;
--		result(18 downto 13) := arg.Eta;
--		result(24 downto 19) := arg.Phi;
--		return result;
--	end function TOB_to_std_logic_vector;

--	function TOB_to_std_logic_vector(arg : JetTOB) return std_logic_vector is
--		variable result : std_logic_vector(19 downto 0);
--	begin
--		--result(18 downto 10) := arg.Et1;
--		result(9 downto 0)   := arg.Et2;
--		result(14 downto 10) := arg.Eta;
--		result(19 downto 15) := arg.Phi;
--		return result;
--	end function TOB_to_std_logic_vector;

--	function TOB_to_std_logic_vector(arg : GenericTOB) return std_logic_vector is
--		variable result : std_logic_vector(21 downto 0);
--	begin
--		result(9 downto 0)   := arg.Et;
--		result(15 downto 10) := arg.eta;
--		result(21 downto 16) := arg.phi;
--		return result;
--	end function TOB_to_std_logic_vector;
	
--	function TOB_to_std_logic_vector(arg : MuonTOB) return std_logic_vector is
--		variable result : std_logic_vector(7 downto 0);
--	begin
--		result(7 downto 5) := arg.Eta;
--		result(4 downto 2) := arg.Phi;
--		result(1 downto 0) := arg.Pt;
--		return result;
--	end function TOB_to_std_logic_vector;

	---------------------------------------------
	-- Functions to convert TOBs to GenericTOB --
	---------------------------------------------
	
	function to_GenericTOB(arg : ClusterTOB) return GenericTOB is
		variable result : GenericTOB;
	begin
		result.Et    := "00" & arg.Et;
		--result.EtSqr := (others => '0');
		result.Eta   := arg.Eta;
		result.Phi   := arg.Phi;
		return result;
	end function to_GenericTOB;
	
	function to_GenericTOB(jet : JetTOB; jet_size : integer) return GenericTOB is
		type JetEtaLut is array (integer range 0 to 31) of integer;
		constant JetEtaTab : JetEtaLut := (
			-39, -- -3.9
			-29, -- -2.95 rounded to -2.9
			-27, -- -2.65 rounded to -2.7
			-25, -- -2.45 rounded to -2.5
			-22, -- -2.2
			-20,
			-18,
			-16,
			-14,
			-12,
			-10,
			-8,
			-6,
			-4,
			-2,
			0,
			2,
			4,
			6,
			8,
			10,
			12,
			14,
			16,
			18,
			20,
			22, -- +2.2
			25, -- +2.45 rounded to 2.5
			27, -- +2.65 rounded to 2.7
			29, -- +2.95 rounded to 2.9
			39, -- +3.9
			39  -- dummy, again +3.9
		);
		variable EtaBin : Integer;
		variable result : GenericTOB;
	begin
		if jet_size = 1 then
			result.Et := '0' & jet.Et1;
		else
			result.Et := jet.Et2;
		end if;
		--result.EtSqr := (others => '0');
		-- convert Eta bins to real eta values
		EtaBin := to_integer(unsigned(jet.Eta));
		result.Eta := std_logic_vector(to_unsigned(JetEtaTab(EtaBin),GenericEtaBitWidth));
		result.Phi   := jet.Phi & '0';
		return result;
	end function to_GenericTOB;

	function to_GenericTOB(arg : MuonTOB) return GenericTOB is --FIXME: Wrong!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
		variable result : GenericTOB;
	begin
		result.Et    := "00000000" & arg.Pt;
		--result.EtSqr := (others => '0');
		result.Eta   := "000" & arg.Eta;
		result.Phi   := "000" & arg.Phi;
		return result;
	end function to_GenericTOB;
	
	function is_in_eta_range(eta_bin : std_logic_vector;
		                      min_bin : std_logic_vector;
		                      max_bin : std_logic_vector) return boolean is
		-- calculate symmetric bin ranges (only needed for forward regions - they are split: low bins and high bins)
		variable eta_max_val : unsigned(eta_bin'length -1 downto 0) := to_unsigned(2**(eta_bin'length) - 1, eta_bin'length);
		variable sym_min_bin : std_logic_vector(eta_bin'length - 1 downto 0) := std_logic_vector(eta_max_val - unsigned(max_bin));
		variable sym_max_bin : std_logic_vector(eta_bin'length - 1 downto 0) := std_logic_vector(eta_max_val - unsigned(min_bin));
		variable result : boolean := false;
	begin
		if ( ((unsigned(eta_bin) >= unsigned(min_bin)) and      -- >= min bin  5bit (32 bins) examples: (0), (14)
		      (unsigned(eta_bin) <= unsigned(max_bin))) or      -- <= max bin                           (5), (17)
		     ((unsigned(eta_bin) >= unsigned(sym_min_bin)) and  -- >= symmetric min bin                (26), (17)
		   	  (unsigned(eta_bin) <= unsigned(sym_max_bin)))     -- <= symmetric max bin                (31), (14)
		   ) then
			result := true;
		else
			result := false;
		end if;
		return result;
	end function is_in_eta_range;

end package body L1TopoFunctions;