-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : gth_quad_multi_gt.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module GTH_QUAD_multi_gt (a Multi GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity GTH_QUAD_multi_gt is
generic
(
    QPLL_FBDIV_TOP                 : integer  := 80;

    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer  := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string   := "FALSE" -- Set to "true" to speed up sim reset
);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    GT0_DRP_BUSY_OUT                        : out  std_logic; 
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt0_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt0_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt0_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt0_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxdlyen_in                          : in   std_logic;
    gt0_rxdlysreset_in                      : in   std_logic;
    gt0_rxdlysresetdone_out                 : out  std_logic;
    gt0_rxphalign_in                        : in   std_logic;
    gt0_rxphaligndone_out                   : out  std_logic;
    gt0_rxphalignen_in                      : in   std_logic;
    gt0_rxphdlyreset_in                     : in   std_logic;
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt0_rxsyncallin_in                      : in   std_logic;
    gt0_rxsyncdone_out                      : out  std_logic;
    gt0_rxsyncin_in                         : in   std_logic;
    gt0_rxsyncmode_in                       : in   std_logic;
    gt0_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt0_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt0_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt0_txdlyen_in                          : in   std_logic;
    gt0_txdlysreset_in                      : in   std_logic;
    gt0_txdlysresetdone_out                 : out  std_logic;
    gt0_txphalign_in                        : in   std_logic;
    gt0_txphaligndone_out                   : out  std_logic;
    gt0_txphalignen_in                      : in   std_logic;
    gt0_txphdlyreset_in                     : in   std_logic;
    gt0_txphinit_in                         : in   std_logic;
    gt0_txphinitdone_out                    : out  std_logic;
    gt0_txsyncallin_in                      : in   std_logic;
    gt0_txsyncdone_out                      : out  std_logic;
    gt0_txsyncin_in                         : in   std_logic;
    gt0_txsyncmode_in                       : in   std_logic;
    gt0_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    GT1_DRP_BUSY_OUT                        : out  std_logic; 
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt1_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt1_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt1_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt1_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxdlyen_in                          : in   std_logic;
    gt1_rxdlysreset_in                      : in   std_logic;
    gt1_rxdlysresetdone_out                 : out  std_logic;
    gt1_rxphalign_in                        : in   std_logic;
    gt1_rxphaligndone_out                   : out  std_logic;
    gt1_rxphalignen_in                      : in   std_logic;
    gt1_rxphdlyreset_in                     : in   std_logic;
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt1_rxsyncallin_in                      : in   std_logic;
    gt1_rxsyncdone_out                      : out  std_logic;
    gt1_rxsyncin_in                         : in   std_logic;
    gt1_rxsyncmode_in                       : in   std_logic;
    gt1_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt1_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt1_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt1_txdlyen_in                          : in   std_logic;
    gt1_txdlysreset_in                      : in   std_logic;
    gt1_txdlysresetdone_out                 : out  std_logic;
    gt1_txphalign_in                        : in   std_logic;
    gt1_txphaligndone_out                   : out  std_logic;
    gt1_txphalignen_in                      : in   std_logic;
    gt1_txphdlyreset_in                     : in   std_logic;
    gt1_txphinit_in                         : in   std_logic;
    gt1_txphinitdone_out                    : out  std_logic;
    gt1_txsyncallin_in                      : in   std_logic;
    gt1_txsyncdone_out                      : out  std_logic;
    gt1_txsyncin_in                         : in   std_logic;
    gt1_txsyncmode_in                       : in   std_logic;
    gt1_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt1_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    GT2_DRP_BUSY_OUT                        : out  std_logic; 
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt2_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt2_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt2_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt2_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxdlyen_in                          : in   std_logic;
    gt2_rxdlysreset_in                      : in   std_logic;
    gt2_rxdlysresetdone_out                 : out  std_logic;
    gt2_rxphalign_in                        : in   std_logic;
    gt2_rxphaligndone_out                   : out  std_logic;
    gt2_rxphalignen_in                      : in   std_logic;
    gt2_rxphdlyreset_in                     : in   std_logic;
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt2_rxsyncallin_in                      : in   std_logic;
    gt2_rxsyncdone_out                      : out  std_logic;
    gt2_rxsyncin_in                         : in   std_logic;
    gt2_rxsyncmode_in                       : in   std_logic;
    gt2_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt2_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt2_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt2_txdlyen_in                          : in   std_logic;
    gt2_txdlysreset_in                      : in   std_logic;
    gt2_txdlysresetdone_out                 : out  std_logic;
    gt2_txphalign_in                        : in   std_logic;
    gt2_txphaligndone_out                   : out  std_logic;
    gt2_txphalignen_in                      : in   std_logic;
    gt2_txphdlyreset_in                     : in   std_logic;
    gt2_txphinit_in                         : in   std_logic;
    gt2_txphinitdone_out                    : out  std_logic;
    gt2_txsyncallin_in                      : in   std_logic;
    gt2_txsyncdone_out                      : out  std_logic;
    gt2_txsyncin_in                         : in   std_logic;
    gt2_txsyncmode_in                       : in   std_logic;
    gt2_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt2_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    GT3_DRP_BUSY_OUT                        : out  std_logic; 
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt3_loopback_in                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    gt3_rxpd_in                             : in   std_logic_vector(1 downto 0);
    gt3_txpd_in                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt3_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxdlyen_in                          : in   std_logic;
    gt3_rxdlysreset_in                      : in   std_logic;
    gt3_rxdlysresetdone_out                 : out  std_logic;
    gt3_rxphalign_in                        : in   std_logic;
    gt3_rxphaligndone_out                   : out  std_logic;
    gt3_rxphalignen_in                      : in   std_logic;
    gt3_rxphdlyreset_in                     : in   std_logic;
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    gt3_rxsyncallin_in                      : in   std_logic;
    gt3_rxsyncdone_out                      : out  std_logic;
    gt3_rxsyncin_in                         : in   std_logic;
    gt3_rxsyncmode_in                       : in   std_logic;
    gt3_rxsyncout_out                       : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt3_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt3_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    gt3_txdlyen_in                          : in   std_logic;
    gt3_txdlysreset_in                      : in   std_logic;
    gt3_txdlysresetdone_out                 : out  std_logic;
    gt3_txphalign_in                        : in   std_logic;
    gt3_txphaligndone_out                   : out  std_logic;
    gt3_txphalignen_in                      : in   std_logic;
    gt3_txphdlyreset_in                     : in   std_logic;
    gt3_txphinit_in                         : in   std_logic;
    gt3_txphinitdone_out                    : out  std_logic;
    gt3_txsyncallin_in                      : in   std_logic;
    gt3_txsyncdone_out                      : out  std_logic;
    gt3_txsyncin_in                         : in   std_logic;
    gt3_txsyncmode_in                       : in   std_logic;
    gt3_txsyncout_out                       : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt3_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);


    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    gt0_gtrefclk0_common_in                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    gt0_qplllock_out                        : out  std_logic;
    gt0_qplllockdetclk_in                   : in   std_logic;
    gt0_qpllpd_in                           : in   std_logic;
    gt0_qpllrefclklost_out                  : out  std_logic;
    gt0_qpllreset_in                        : in   std_logic


);


end GTH_QUAD_multi_gt;
    
architecture RTL of GTH_QUAD_multi_gt is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "GTH_QUAD_multi_gt,gtwizard_v2_6,{protocol_file=Start_from_scratch}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
signal  tied_to_ground_i                :   std_logic;
signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
signal  tied_to_vcc_i                   :   std_logic;
signal   gt0_qplloutclk_i         :   std_logic;
signal   gt0_qplloutrefclk_i      :   std_logic;

signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
 

signal   gt0_qpllclk_i            :   std_logic;
signal   gt0_qpllrefclk_i         :   std_logic;
    signal    gt0_rst_i                       : std_logic;
signal   gt1_qpllclk_i            :   std_logic;
signal   gt1_qpllrefclk_i         :   std_logic;
    signal    gt1_rst_i                       : std_logic;
signal   gt2_qpllclk_i            :   std_logic;
signal   gt2_qpllrefclk_i         :   std_logic;
    signal    gt2_rst_i                       : std_logic;
signal   gt3_qpllclk_i            :   std_logic;
signal   gt3_qpllrefclk_i         :   std_logic;
    signal    gt3_rst_i                       : std_logic;


--*************************** Component Declarations **************************
component GTH_QUAD_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP    : string := "FALSE";
    EXAMPLE_SIMULATION        : integer  := 0;   
    TXSYNC_OVRD_IN            : bit    := '0';
    TXSYNC_MULTILANE_IN       : bit    := '0'     
);
port 
(   
    RST_IN                                  : in   std_logic;
    DRP_BUSY_OUT                            : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    drpaddr_in                              : in   std_logic_vector(8 downto 0);
    drpclk_in                               : in   std_logic;
    drpdi_in                                : in   std_logic_vector(15 downto 0);
    drpdo_out                               : out  std_logic_vector(15 downto 0);
    drpen_in                                : in   std_logic;
    drprdy_out                              : out  std_logic;
    drpwe_in                                : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    qpllclk_in                              : in   std_logic;
    qpllrefclk_in                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    loopback_in                             : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    rxpd_in                                 : in   std_logic_vector(1 downto 0);
    txpd_in                                 : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    rxuserrdy_in                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    eyescandataerror_out                    : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    rxcdrlock_out                           : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    rxusrclk_in                             : in   std_logic;
    rxusrclk2_in                            : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    rxdata_out                              : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    rxdisperr_out                           : out  std_logic_vector(3 downto 0);
    rxnotintable_out                        : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gthrxn_in                               : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    rxdlyen_in                              : in   std_logic;
    rxdlysreset_in                          : in   std_logic;
    rxdlysresetdone_out                     : out  std_logic;
    rxphalign_in                            : in   std_logic;
    rxphaligndone_out                       : out  std_logic;
    rxphalignen_in                          : in   std_logic;
    rxphdlyreset_in                         : in   std_logic;
    rxphmonitor_out                         : out  std_logic_vector(4 downto 0);
    rxphslipmonitor_out                     : out  std_logic_vector(4 downto 0);
    rxsyncallin_in                          : in   std_logic;
    rxsyncdone_out                          : out  std_logic;
    rxsyncin_in                             : in   std_logic;
    rxsyncmode_in                           : in   std_logic;
    rxsyncout_out                           : out  std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    rxmcommaalignen_in                      : in   std_logic;
    rxpcommaalignen_in                      : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    rxlpmhfhold_in                          : in   std_logic;
    rxlpmlfhold_in                          : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    rxoutclk_out                            : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gtrxreset_in                            : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    rxcharisk_out                           : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gthrxp_in                               : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    rxresetdone_out                         : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    txpostcursor_in                         : in   std_logic_vector(4 downto 0);
    txprecursor_in                          : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gttxreset_in                            : in   std_logic;
    txuserrdy_in                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    txusrclk_in                             : in   std_logic;
    txusrclk2_in                            : in   std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    txdlyen_in                              : in   std_logic;
    txdlysreset_in                          : in   std_logic;
    txdlysresetdone_out                     : out  std_logic;
    txphalign_in                            : in   std_logic;
    txphaligndone_out                       : out  std_logic;
    txphalignen_in                          : in   std_logic;
    txphdlyreset_in                         : in   std_logic;
    txphinit_in                             : in   std_logic;
    txphinitdone_out                        : out  std_logic;
    txsyncallin_in                          : in   std_logic;
    txsyncdone_out                          : out  std_logic;
    txsyncin_in                             : in   std_logic;
    txsyncmode_in                           : in   std_logic;
    txsyncout_out                           : out  std_logic;
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    txdiffctrl_in                           : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    txdata_in                               : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gthtxn_out                              : out  std_logic;
    gthtxp_out                              : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    txoutclk_out                            : out  std_logic;
    txoutclkfabric_out                      : out  std_logic;
    txoutclkpcs_out                         : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    txresetdone_out                         : out  std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    txcharisk_in                            : in   std_logic_vector(3 downto 0)


);
end component;


--*************************Logic to set Attribute QPLL_FB_DIV*****************************
    impure function conv_qpll_fbdiv_top (qpllfbdiv_top : in integer) return bit_vector is
    begin
       if (qpllfbdiv_top = 16) then
         return "0000100000";
       elsif (qpllfbdiv_top = 20) then
         return "0000110000" ;
       elsif (qpllfbdiv_top = 32) then
         return "0001100000" ;
       elsif (qpllfbdiv_top = 40) then
         return "0010000000" ;
       elsif (qpllfbdiv_top = 64) then
         return "0011100000" ;
       elsif (qpllfbdiv_top = 66) then
         return "0101000000" ;
       elsif (qpllfbdiv_top = 80) then
         return "0100100000" ;
       elsif (qpllfbdiv_top = 100) then
         return "0101110000" ;
       else 
         return "0000000000" ;
       end if;
    end function;

    impure function conv_qpll_fbdiv_ratio (qpllfbdiv_top : in integer) return bit is
    begin
       if (qpllfbdiv_top = 16) then
         return '1';
       elsif (qpllfbdiv_top = 20) then
         return '1' ;
       elsif (qpllfbdiv_top = 32) then
         return '1' ;
       elsif (qpllfbdiv_top = 40) then
         return '1' ;
       elsif (qpllfbdiv_top = 64) then
         return '1' ;
       elsif (qpllfbdiv_top = 66) then
         return '0' ;
       elsif (qpllfbdiv_top = 80) then
         return '1' ;
       elsif (qpllfbdiv_top = 100) then
         return '1' ;
       else 
         return '1' ;
       end if;
    end function;

    constant   QPLL_FBDIV_IN    :   bit_vector(9 downto 0) := conv_qpll_fbdiv_top(QPLL_FBDIV_TOP);
    constant   QPLL_FBDIV_RATIO :   bit := conv_qpll_fbdiv_ratio(QPLL_FBDIV_TOP);

--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_qpllclk_i    <= gt0_qplloutclk_i;  
    gt0_qpllrefclk_i <= gt0_qplloutrefclk_i; 
    gt1_qpllclk_i    <= gt0_qplloutclk_i;  
    gt1_qpllrefclk_i <= gt0_qplloutrefclk_i; 
    gt2_qpllclk_i    <= gt0_qplloutclk_i;  
    gt2_qpllrefclk_i <= gt0_qplloutrefclk_i; 
    gt3_qpllclk_i    <= gt0_qplloutclk_i;  
    gt3_qpllrefclk_i <= gt0_qplloutrefclk_i; 

      gt0_rst_i        <= GT0_QPLLRESET_IN;
   
      gt1_rst_i        <= GT0_QPLLRESET_IN;
   
      gt2_rst_i        <= GT0_QPLLRESET_IN;
   
      gt3_rst_i        <= GT0_QPLLRESET_IN;
   
     

    --------------------------- GT Instances  -------------------------------   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
gt0_GTH_QUAD_i : GTH_QUAD_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt0_rst_i,
        DRP_BUSY_OUT                    =>      GT0_DRP_BUSY_OUT,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt0_drpaddr_in,
        drpclk_in                       =>      gt0_drpclk_in,
        drpdi_in                        =>      gt0_drpdi_in,
        drpdo_out                       =>      gt0_drpdo_out,
        drpen_in                        =>      gt0_drpen_in,
        drprdy_out                      =>      gt0_drprdy_out,
        drpwe_in                        =>      gt0_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt0_qpllclk_i,
        qpllrefclk_in                   =>      gt0_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        loopback_in                     =>      gt0_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        rxpd_in                         =>      gt0_rxpd_in,
        txpd_in                         =>      gt0_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        rxuserrdy_in                    =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt0_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        rxcdrlock_out                   =>      gt0_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt0_rxusrclk_in,
        rxusrclk2_in                    =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt0_rxdisperr_out,
        rxnotintable_out                =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt0_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt0_rxdlyen_in,
        rxdlysreset_in                  =>      gt0_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt0_rxdlysresetdone_out,
        rxphalign_in                    =>      gt0_rxphalign_in,
        rxphaligndone_out               =>      gt0_rxphaligndone_out,
        rxphalignen_in                  =>      gt0_rxphalignen_in,
        rxphdlyreset_in                 =>      gt0_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt0_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt0_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt0_rxsyncallin_in,
        rxsyncdone_out                  =>      gt0_rxsyncdone_out,
        rxsyncin_in                     =>      gt0_rxsyncin_in,
        rxsyncmode_in                   =>      gt0_rxsyncmode_in,
        rxsyncout_out                   =>      gt0_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxmcommaalignen_in              =>      gt0_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt0_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt0_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt0_rxlpmlfhold_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt0_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt0_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt0_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt0_rxresetdone_out,
        ------------------------ TX Configurable Driver Ports ----------------------
        txpostcursor_in                 =>      gt0_txpostcursor_in,
        txprecursor_in                  =>      gt0_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt0_gttxreset_in,
        txuserrdy_in                    =>      gt0_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt0_txusrclk_in,
        txusrclk2_in                    =>      gt0_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt0_txdlyen_in,
        txdlysreset_in                  =>      gt0_txdlysreset_in,
        txdlysresetdone_out             =>      gt0_txdlysresetdone_out,
        txphalign_in                    =>      gt0_txphalign_in,
        txphaligndone_out               =>      gt0_txphaligndone_out,
        txphalignen_in                  =>      gt0_txphalignen_in,
        txphdlyreset_in                 =>      gt0_txphdlyreset_in,
        txphinit_in                     =>      gt0_txphinit_in,
        txphinitdone_out                =>      gt0_txphinitdone_out,
        txsyncallin_in                  =>      gt0_txsyncallin_in,
        txsyncdone_out                  =>      gt0_txsyncdone_out,
        txsyncin_in                     =>      gt0_txsyncin_in,
        txsyncmode_in                   =>      gt0_txsyncmode_in,
        txsyncout_out                   =>      gt0_txsyncout_out,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        txdiffctrl_in                   =>      gt0_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt0_gthtxn_out,
        gthtxp_out                      =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt0_txoutclk_out,
        txoutclkfabric_out              =>      gt0_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt0_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt0_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y1)
gt1_GTH_QUAD_i : GTH_QUAD_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt1_rst_i,
        DRP_BUSY_OUT                    =>      GT1_DRP_BUSY_OUT,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt1_drpaddr_in,
        drpclk_in                       =>      gt1_drpclk_in,
        drpdi_in                        =>      gt1_drpdi_in,
        drpdo_out                       =>      gt1_drpdo_out,
        drpen_in                        =>      gt1_drpen_in,
        drprdy_out                      =>      gt1_drprdy_out,
        drpwe_in                        =>      gt1_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt1_qpllclk_i,
        qpllrefclk_in                   =>      gt1_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        loopback_in                     =>      gt1_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        rxpd_in                         =>      gt1_rxpd_in,
        txpd_in                         =>      gt1_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        rxuserrdy_in                    =>      gt1_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt1_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        rxcdrlock_out                   =>      gt1_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt1_rxusrclk_in,
        rxusrclk2_in                    =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt1_rxdisperr_out,
        rxnotintable_out                =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt1_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt1_rxdlyen_in,
        rxdlysreset_in                  =>      gt1_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt1_rxdlysresetdone_out,
        rxphalign_in                    =>      gt1_rxphalign_in,
        rxphaligndone_out               =>      gt1_rxphaligndone_out,
        rxphalignen_in                  =>      gt1_rxphalignen_in,
        rxphdlyreset_in                 =>      gt1_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt1_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt1_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt1_rxsyncallin_in,
        rxsyncdone_out                  =>      gt1_rxsyncdone_out,
        rxsyncin_in                     =>      gt1_rxsyncin_in,
        rxsyncmode_in                   =>      gt1_rxsyncmode_in,
        rxsyncout_out                   =>      gt1_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxmcommaalignen_in              =>      gt1_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt1_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt1_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt1_rxlpmlfhold_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt1_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt1_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt1_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt1_rxresetdone_out,
        ------------------------ TX Configurable Driver Ports ----------------------
        txpostcursor_in                 =>      gt1_txpostcursor_in,
        txprecursor_in                  =>      gt1_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt1_gttxreset_in,
        txuserrdy_in                    =>      gt1_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt1_txusrclk_in,
        txusrclk2_in                    =>      gt1_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt1_txdlyen_in,
        txdlysreset_in                  =>      gt1_txdlysreset_in,
        txdlysresetdone_out             =>      gt1_txdlysresetdone_out,
        txphalign_in                    =>      gt1_txphalign_in,
        txphaligndone_out               =>      gt1_txphaligndone_out,
        txphalignen_in                  =>      gt1_txphalignen_in,
        txphdlyreset_in                 =>      gt1_txphdlyreset_in,
        txphinit_in                     =>      gt1_txphinit_in,
        txphinitdone_out                =>      gt1_txphinitdone_out,
        txsyncallin_in                  =>      gt1_txsyncallin_in,
        txsyncdone_out                  =>      gt1_txsyncdone_out,
        txsyncin_in                     =>      gt1_txsyncin_in,
        txsyncmode_in                   =>      gt1_txsyncmode_in,
        txsyncout_out                   =>      gt1_txsyncout_out,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        txdiffctrl_in                   =>      gt1_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt1_gthtxn_out,
        gthtxp_out                      =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt1_txoutclk_out,
        txoutclkfabric_out              =>      gt1_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt1_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt1_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt1_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y2)
gt2_GTH_QUAD_i : GTH_QUAD_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt2_rst_i,
        DRP_BUSY_OUT                    =>      GT2_DRP_BUSY_OUT,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt2_drpaddr_in,
        drpclk_in                       =>      gt2_drpclk_in,
        drpdi_in                        =>      gt2_drpdi_in,
        drpdo_out                       =>      gt2_drpdo_out,
        drpen_in                        =>      gt2_drpen_in,
        drprdy_out                      =>      gt2_drprdy_out,
        drpwe_in                        =>      gt2_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt2_qpllclk_i,
        qpllrefclk_in                   =>      gt2_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        loopback_in                     =>      gt2_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        rxpd_in                         =>      gt2_rxpd_in,
        txpd_in                         =>      gt2_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        rxuserrdy_in                    =>      gt2_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt2_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        rxcdrlock_out                   =>      gt2_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt2_rxusrclk_in,
        rxusrclk2_in                    =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt2_rxdisperr_out,
        rxnotintable_out                =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt2_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt2_rxdlyen_in,
        rxdlysreset_in                  =>      gt2_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt2_rxdlysresetdone_out,
        rxphalign_in                    =>      gt2_rxphalign_in,
        rxphaligndone_out               =>      gt2_rxphaligndone_out,
        rxphalignen_in                  =>      gt2_rxphalignen_in,
        rxphdlyreset_in                 =>      gt2_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt2_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt2_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt2_rxsyncallin_in,
        rxsyncdone_out                  =>      gt2_rxsyncdone_out,
        rxsyncin_in                     =>      gt2_rxsyncin_in,
        rxsyncmode_in                   =>      gt2_rxsyncmode_in,
        rxsyncout_out                   =>      gt2_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxmcommaalignen_in              =>      gt2_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt2_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt2_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt2_rxlpmlfhold_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt2_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt2_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt2_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt2_rxresetdone_out,
        ------------------------ TX Configurable Driver Ports ----------------------
        txpostcursor_in                 =>      gt2_txpostcursor_in,
        txprecursor_in                  =>      gt2_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt2_gttxreset_in,
        txuserrdy_in                    =>      gt2_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt2_txusrclk_in,
        txusrclk2_in                    =>      gt2_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt2_txdlyen_in,
        txdlysreset_in                  =>      gt2_txdlysreset_in,
        txdlysresetdone_out             =>      gt2_txdlysresetdone_out,
        txphalign_in                    =>      gt2_txphalign_in,
        txphaligndone_out               =>      gt2_txphaligndone_out,
        txphalignen_in                  =>      gt2_txphalignen_in,
        txphdlyreset_in                 =>      gt2_txphdlyreset_in,
        txphinit_in                     =>      gt2_txphinit_in,
        txphinitdone_out                =>      gt2_txphinitdone_out,
        txsyncallin_in                  =>      gt2_txsyncallin_in,
        txsyncdone_out                  =>      gt2_txsyncdone_out,
        txsyncin_in                     =>      gt2_txsyncin_in,
        txsyncmode_in                   =>      gt2_txsyncmode_in,
        txsyncout_out                   =>      gt2_txsyncout_out,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        txdiffctrl_in                   =>      gt2_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt2_gthtxn_out,
        gthtxp_out                      =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt2_txoutclk_out,
        txoutclkfabric_out              =>      gt2_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt2_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt2_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt2_txcharisk_in

    );
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y3)
gt3_GTH_QUAD_i : GTH_QUAD_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('1'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt3_rst_i,
        DRP_BUSY_OUT                    =>      GT3_DRP_BUSY_OUT,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt3_drpaddr_in,
        drpclk_in                       =>      gt3_drpclk_in,
        drpdi_in                        =>      gt3_drpdi_in,
        drpdo_out                       =>      gt3_drpdo_out,
        drpen_in                        =>      gt3_drpen_in,
        drprdy_out                      =>      gt3_drprdy_out,
        drpwe_in                        =>      gt3_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt3_qpllclk_i,
        qpllrefclk_in                   =>      gt3_qpllrefclk_i,
        ------------------------------- Loopback Ports -----------------------------
        loopback_in                     =>      gt3_loopback_in,
        ------------------------------ Power-Down Ports ----------------------------
        rxpd_in                         =>      gt3_rxpd_in,
        txpd_in                         =>      gt3_txpd_in,
        --------------------- RX Initialization and Reset Ports --------------------
        rxuserrdy_in                    =>      gt3_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt3_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        rxcdrlock_out                   =>      gt3_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt3_rxusrclk_in,
        rxusrclk2_in                    =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt3_rxdisperr_out,
        rxnotintable_out                =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt3_gthrxn_in,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        rxdlyen_in                      =>      gt3_rxdlyen_in,
        rxdlysreset_in                  =>      gt3_rxdlysreset_in,
        rxdlysresetdone_out             =>      gt3_rxdlysresetdone_out,
        rxphalign_in                    =>      gt3_rxphalign_in,
        rxphaligndone_out               =>      gt3_rxphaligndone_out,
        rxphalignen_in                  =>      gt3_rxphalignen_in,
        rxphdlyreset_in                 =>      gt3_rxphdlyreset_in,
        rxphmonitor_out                 =>      gt3_rxphmonitor_out,
        rxphslipmonitor_out             =>      gt3_rxphslipmonitor_out,
        rxsyncallin_in                  =>      gt3_rxsyncallin_in,
        rxsyncdone_out                  =>      gt3_rxsyncdone_out,
        rxsyncin_in                     =>      gt3_rxsyncin_in,
        rxsyncmode_in                   =>      gt3_rxsyncmode_in,
        rxsyncout_out                   =>      gt3_rxsyncout_out,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxmcommaalignen_in              =>      gt3_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt3_rxpcommaalignen_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt3_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt3_rxlpmlfhold_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt3_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt3_gtrxreset_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt3_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt3_rxresetdone_out,
        ------------------------ TX Configurable Driver Ports ----------------------
        txpostcursor_in                 =>      gt3_txpostcursor_in,
        txprecursor_in                  =>      gt3_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt3_gttxreset_in,
        txuserrdy_in                    =>      gt3_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt3_txusrclk_in,
        txusrclk2_in                    =>      gt3_txusrclk2_in,
        ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
        txdlyen_in                      =>      gt3_txdlyen_in,
        txdlysreset_in                  =>      gt3_txdlysreset_in,
        txdlysresetdone_out             =>      gt3_txdlysresetdone_out,
        txphalign_in                    =>      gt3_txphalign_in,
        txphaligndone_out               =>      gt3_txphaligndone_out,
        txphalignen_in                  =>      gt3_txphalignen_in,
        txphdlyreset_in                 =>      gt3_txphdlyreset_in,
        txphinit_in                     =>      gt3_txphinit_in,
        txphinitdone_out                =>      gt3_txphinitdone_out,
        txsyncallin_in                  =>      gt3_txsyncallin_in,
        txsyncdone_out                  =>      gt3_txsyncdone_out,
        txsyncin_in                     =>      gt3_txsyncin_in,
        txsyncmode_in                   =>      gt3_txsyncmode_in,
        txsyncout_out                   =>      gt3_txsyncout_out,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        txdiffctrl_in                   =>      gt3_txdiffctrl_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt3_gthtxn_out,
        gthtxp_out                      =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt3_txoutclk_out,
        txoutclkfabric_out              =>      gt3_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt3_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt3_txresetdone_out,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt3_txcharisk_in

    );
    

    --_________________________________________________________________________
    --_________________________________________________________________________
    --_________________________GTHE2_COMMON____________________________________

    gthe2_common_0_i : GTHE2_COMMON
    generic map
    (
            -- Simulation attributes
            SIM_RESET_SPEEDUP    => WRAPPER_SIM_GTRESET_SPEEDUP,
            SIM_QPLLREFCLK_SEL   => ("001"),
            SIM_VERSION          => ("2.0"),


       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000040000001050"),
        COMMON_CFG                              =>     (x"00000000"),
        QPLL_CFG                                =>     (x"04801C7"),
        QPLL_CLKOUT_CFG                         =>     ("1111"),
        QPLL_COARSE_FREQ_OVRD                   =>     ("010000"),
        QPLL_COARSE_FREQ_OVRD_EN                =>     ('0'),
        QPLL_CP                                 =>     ("0000011111"),
        QPLL_CP_MONITOR_EN                      =>     ('0'),
        QPLL_DMONITOR_SEL                       =>     ('0'),
        QPLL_FBDIV                              =>     (QPLL_FBDIV_IN),
        QPLL_FBDIV_MONITOR_EN                   =>     ('0'),
        QPLL_FBDIV_RATIO                        =>     (QPLL_FBDIV_RATIO),
        QPLL_INIT_CFG                           =>     (x"000006"),
        QPLL_LOCK_CFG                           =>     (x"05E8"),
        QPLL_LPF                                =>     ("1111"),
        QPLL_REFCLK_DIV                         =>     (1),
        RSVD_ATTR0                              =>     (x"0000"),
        RSVD_ATTR1                              =>     (x"0000"),
        QPLL_RP_COMP                            =>     ('0'),
        QPLL_VTRL_RESET                         =>     ("00"),
        RCAL_CFG                                =>     ("00")

        
    )
    port map
    (
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GTGREFCLK                       =>      tied_to_ground_i,
        GTNORTHREFCLK0                  =>      tied_to_ground_i,
        GTNORTHREFCLK1                  =>      tied_to_ground_i,
        GTREFCLK0                       =>      gt0_gtrefclk0_common_in,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTSOUTHREFCLK0                  =>      tied_to_ground_i,
        GTSOUTHREFCLK1                  =>      tied_to_ground_i,
        ------------------------- Common Block -  QPLL Ports -----------------------
        QPLLDMONITOR                    =>      open,
        ----------------------- Common Block - Clocking Ports ----------------------
        QPLLOUTCLK                      =>      gt0_qplloutclk_i,
        QPLLOUTREFCLK                   =>      gt0_qplloutrefclk_i,
        REFCLKOUTMONITOR                =>      open,
        ------------------------- Common Block - QPLL Ports ------------------------
        BGRCALOVRDENB                   =>      tied_to_vcc_i,
        PMARSVDOUT                      =>      open,
        QPLLFBCLKLOST                   =>      open,
        QPLLLOCK                        =>      gt0_qplllock_out,
        QPLLLOCKDETCLK                  =>      gt0_qplllockdetclk_in,
        QPLLLOCKEN                      =>      tied_to_vcc_i,
        QPLLOUTRESET                    =>      tied_to_ground_i,
        QPLLPD                          =>      gt0_qpllpd_in,
        QPLLREFCLKLOST                  =>      gt0_qpllrefclklost_out,
        QPLLREFCLKSEL                   =>      "001",
        QPLLRESET                       =>      gt0_qpllreset_in,
        QPLLRSVD1                       =>      "0000000000000000",
        QPLLRSVD2                       =>      "11111",
        --------------------------------- QPLL Ports -------------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i

    );

end RTL;
     
