-------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : gtx_quad_no_buffer_config_gtmodel.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gtx_quad_no_buffer_config_gtmodel 
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 

-- Use this file for fast simulation mode setup                              
-------------------------------------------------------------------------------
library unisim;
library unifast;

configuration gtx_quad_no_buffer_TB_cfg of gtx_quad_no_buffer_TB is
for RTL
  for gtx_quad_no_buffer_exdes_i:gtx_quad_no_buffer_exdes
    use entity work.gtx_quad_no_buffer_exdes;
    for RTL
       for gtx_quad_no_buffer_init_i:gtx_quad_no_buffer_init
          use entity work.gtx_quad_no_buffer_init;
          for RTL
             for gtx_quad_no_buffer_i:gtx_quad_no_buffer
                use entity work.gtx_quad_no_buffer;
                for RTL
                   for gt0_gtx_quad_no_buffer_i:gtx_quad_no_buffer_GT
                      use entity work.gtx_quad_no_buffer_GT;
                      for RTL
                          for all:GTXE2_CHANNEL
                             use entity unifast.GTXE2_CHANNEL;
                          end for;
                      end for;
                   end for;
                end for;
             end for;
          end for;
       end for;
    end for;
  end for;
end for;
end gtx_quad_no_buffer_TB_cfg;

