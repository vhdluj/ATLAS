`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Iu14w2w0KSVQJh5kTz2fDmW/Yq777xPAuiY1c9H5g4XbHzVHRC97+NicvtifFQDa2iFSXBVGYhf9
oMWIWKga+w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jWn20MlwOXOCSfHGQ4KhVv2t9i6tMMYIF66b6nc/0DsIWgkn1DIpVa8KX6lfxU9RFEfRGHgpBJAS
JUTGqFBS9CFePmeSvnzrRnyQVGcTDNNizbPbNMoBZOLQTHnPJuBgise7lbYAZ3mbWpLrl7/0fGhp
EwHdoKU2SVtPIljp+4o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nelQ8WUHWgZ9dCdDGLoD10m+XhgDJfyZCRdMfuOyeBhjpMBZV/oGL3neCSJzXOwn178Lqeryzf8+
aIcaSF9A36X0NO240hWXTuee0ZP/0BEFoV1uIJBUDffP0kL48Bhc0L1IGjIZdu/z/J5DgljV5wPf
QFbf+stAsADdUSbWvlaerhL1cqRT7a5TmSGUO+9M0u9qV8hiuzkSDOT5OZXCqCJbDoeS4oZvWJ/I
K/ZmE9pdeQCtbzLK7Q9VuWbsLid8qL33pge7eMZnv6cgZTGIb7PTUrJdcRU6+P2MW+JDvJh+x5WS
rDpuu0AHaDR6wo/ol6/0PEj7TW/yj03beTQqBg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hXF4yyX6GXXJbUfC9ZzCVwLmcNrSoizKfnMaaXAHTexx0tk+FAOXPobEfBLpySdSYv+n82Ivg5EA
vvVmkRFX4WbnZxGJ5cGPgBehv0Ecw9fWzoE3NyK87Uo7Tx2nF2TBcpQqd+mDt1hZc22inNFSMEro
rfctizRxfnHdHUzkqSo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hEVvwe7AIuj2L7eQYfxXyNUwo0dzWKYwCHfe6lsxFgtMvVQnpjkc6AsbsVSG+mhR3lMUMUuQD/H4
VZqTY/PNksrpZW2XNUbqVXvWKMWRLbXzlsE3E0wZp1cOD+sCi3oa7d5/eqK5/Ew60cfchCt4XMFX
p1/wBNaxZr6/wnQNIjyBt/L1AGsnuu6DwMje7ZUuw+rFt5g7y8PZEbi+rEHsCQUeA7c0SFBlUfsE
b7HNrDU3s/Sqi5//4gZNX1AcGEg9ReJh+7hbqbDaqs43tqBDW87Cvz7VrqgMkqsGYdr5+D1fk8Lp
I4pxZ4tcMa8J3A9YNqwQY92RjdVMhBuDbJK44Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19568)
`protect data_block
iTN29yBmNSKMHd6B7/cU8wojIl/aWOTapYfXWsS3837v++RJ2IgzyAjq3/AerEP2/8N1I8QLJiD4
RFpzzSIuMJkC7QJOFzTdW/hOPms8e4HItD0fNAs4gmWrJIzYahJH0Sdi/s0HA0AiLWnrhjFPMLos
FmObTpehMS8ldunSXA7Hf4bIgK00JUfMoVDHZxaBnj8qDkxfz2qACbPDGvOwco71zsoeZpoPJXPA
GKogA3be7DaA79FMeB8XKDlW4PONvUvW9uadSuX8E4GxtfEixy1rL4yUchb9kGQKa5f2WIuQXmi9
xyVQsxtiM3waKLHEBEcoj43Pj7Q2NCcnv2DVJeHg57b2iO2uvH/6aQgbYOTyxYnD4zAOoHHFNXCC
yt90HnawvWemAEEeD/8OpEiiUxRBY+xW+r4qs1XUSeJmNNxSN+BFIw0I36os24c4AMFgpmjlxgYv
pfLBpuk23CDgFspwvKYhsT+9jIWp98m15FUHwXr5rcs8SItdw6p+jmo4sAN/7clQUghodF/VyNuD
w0Ls+eSeXqhxu8zeUgdJkPPek4enCy1fnAgfok/65HdgiEWd2c9d7g6luj9jWPawcqqkDKbgoBBs
91fIZJkG77yB+jJ70/Ct4pDtB0SJelVibR7BY0r+ZvR/PakURR9N6Qhv/rqiXLAXTVSkXWjknonV
bZ2wIS37pzcaX1cQeFzudZLHG/n4nlA1nn6UvdCx7iIYxm8+0r9OyhZ00mpvbj2sjGXIltHDfaAm
VKe1yBEMTanhjF/w0mdkUcBq77jUb4+T/Dm4H+ODcxL3VYxh4fquiudY6o/ovSLfhzXg9o5f1QWX
us/lImAgxRACwyr6obdwxnebth1YmOFOyi8gkvDlqexZNFnirTmumyPyDzWXX9p52UZvn4i1oQPL
QFNkgCN431BzCgO8YONBZ353tuaaFOoFqfySo5Sgrwjfd0yhF1+wGMzBFkJ15OYkSq1SCZMzH1IP
AHHsclYOlxC9IJcMiPEUWspE4kgIiaKQ0k1k6yH/2Ze7ph1BuENAQjJlRl75w1nGOinKKAkh5W+h
bK7Et8ITYHGxjENg6zQKw+NNXVN3XqjmVgS/lNdkaysaqvCJOisbTL/6iXQDf4jNm7VvLfqpZLHT
EZdbvv8zD35sz8lbvkPdrWz1tEstFyyEtTCRULL6KFZcdX1pWGBWQIxURd7YBzKyI5jW3m9z5xra
SszgBsA3KimWuUwspVdFcZwiY9Xur9H5xkZ/qU/z141xa1wEQ2QYs0094pzpwSk7ePwuIld86dU3
iHkvTtneoPwj8oqGKViLcvWu+r7+GCJlJCHrSugDflf1pfEgL7yJ8r+7sfmjUlb9fvAwFi5ilNnN
fZCeJw1rwZ/uFP3zAD467A2OCvgg0gU3Z69aEWWYuiR+NN3ciR822zioN+qJjC/3qgsQNfuOTsmA
eyFB5wzJZ8/BEOwHz/1jNfUcHHN9NuBADM/EePM2RCylypjK+upz13TBMzp2ikkg0HfUDjSwLnGC
QHo2zkgYDTqE/7yN2Gffu4qhrM1Ck4123k+nOKFgCkt8/OwSRjM2+9vla9z/+eN8kTyLoWTeA5p2
ucKhbcIau/0Ne36QVW9REaujTCmkq+TZJSZXa5AoDSCTbDc+NKJpO+7T7xE2V/CUAqaq9eflyEA/
hpRynFXjq0Cg6Lfj0yP8BpvnIIpKas3kzlrGzksc9vrVnYQE2BpQKHBckHGDP3jS4YedwsCo9ONx
4VU2XPX+bayWy3JqZRm37KomS24NtFwCtNTKyz0PFdmdkLSFjnoH5RaWBgzSYO/D/Z9Q6c+rd7jh
DT8x9ZnkiYvlxJC3QAP2RODqyIBMZz+aQZW8eX/Eq4t1iJKzF+QVqIH0ejWuGsMRg4GXtEHA9lqV
JErKiPgjEwZuK0tAI29MdrQlOOIsd3RVFZ4VekUtFDDYZyR/bqwI0H2t+/krRbDqbETK2WYLACRv
ohFF7kDwJ92ES8HrMbQFAgnU1RLQiSRr3ILrEacRpDipAhhIsK53ZEERXMH1e2uLk+NgkcWGEklO
vA8qhJWLmYzC46OFlMfGudiygIX7g38j1AVeBSbrmAQF5P3g/HXdaJjJMWyRnst3cmkRtw0Zb1Ch
mG+/AJMEHClGqKpHizoQeCIQkppnx/5faf7+I9jCgIbSLh7L3HRZ6TcqvhUSR+qvCi8sF93eEbd4
IueXl5h9qbn9Dnk4JUw+NDE73kA+0BVLQ/i0Rxct/WkDoZBc9Ym8pA/3fGUTJT0BVdnY8HiOmnaq
uBcQf4UVhuTjctjYg4NzkpAl29E+FYZoX2oqWqu43PQhRkLYDGzqBDPK04BV2MZhvn9vGZZRlceB
d1JD2ma6mzJi4alAN+ZBkl+81ZkMygD5A+HZt3jXlPMkEyx3agc0KJYXCoAslp0pi00fpmQWFmBn
k1PTWjuh5/BWlHAtoI1zYmLFL3OwsgfdVj6Usmtmif1kkgc9SQiz+/RnXfxuXSm2LC6SgnEGiohz
izY1DqL+RvdNJGBE1W6G994VUGlD7IfDTENT8D0FktenG0YLBhgyb9rbWbqDtP/GVxyqcEBHJmft
axtOpNNvIBZwV/ms4U7KVGMfv/AZR+YjVzqe6M1eXeGhwyvAwIz2w1aa7yTWvVYTeJOvCkHYhrd0
uQrwHq+dXikDi8gRlt/MWI+E0HUPBdr+5Kxo5N1wannXEIW0+PvNGxvw5j7dBEI/JE5WgZk1AJsm
iTsEgVuA56qKw5VHj7+E0GRhz3v/1sArkN0QXC2+imMxamq0qwhg8xzVolFMYsZgO48eSTUvgMmC
+5abkG0ewy/dCKDd3KPyqi0flNY+9hp81r0wE7AQDUim032VekvVlwec+LfZWWP/iPu1UMLg5N16
kaQHS4vypeNPftK68fw9oG6zJ2cs9aJ/UCE7OcCu1lVe/iJuvzJ9u7dXCmVaD0wI/BaGq5wnd0Eb
DEQIKcYnR59bqO+NJm4jaJCLuANowUHcx9fLy/9NAUMILeqe6EE4hv4Rt3+Nm1uD0GkNvrYA0aEa
Nu8IcmGFdkIRKLOub7EiqWLs26caunn4OCTbNqmBAUwr1RkiHPJvMhf77t5gdC1zmYPU2xJ05j+z
VhBsE81HBshPGDXQoemlhdgYXnDkwwfYIohPOpQSAUOw/k+yV7JlmAFD6wZ7f2cJLLgHqQ0Zr6VD
Pi6fTaAFOvNw9RMFnoZ9OBxTPZEcQuGhX0+Fm53gXbteRdNFhihAEPzVftvNTjD9n7Z7+yyHxUf3
MNWCbcYQka/QmQwM0Uq9NbYLjjt3dkZcFW2o78Q5ChAjSbD+ERH7ujOn7/JwmKql4kyfhop50s09
kRWKrEe31UYKmHcDLKMdDnH6VPZl4p0Zq6hQnKXqwc/JxWhbJWDC216jg/CLC1SShlNK56Uf4Xb+
i8PxmRCvnh7+GVEsqohtlkZDl35C09ae2QHdUVg2C9qsrTB4lQqNoVFZOugd+xZ9f9A4GrTl/t2Z
dlQxeeE9kahw3ZX+CpjJeb77JD4tbKMIxJoOi4nB02t1k6V7PXAhri7yRMsr7mtm6/kNEANKxNNU
OgRAbaI/CMXjC/yE123U+9ioton3uMUn4AXPe8dJeRz/m/boivtlNYV/7j3t+PGDAyCcTKZW21me
iARY6jY5pnpK1xYwhcyLWCSJteBrkdDkPs7dXVf6sxdbY+zkW7nkHqe664hxo06kU0tvfZoOHkXD
O8g26pUtbjI7RSt+Yuh6T2PCP/p+D6a/uqoW6XFkf68Y9NHTnetC+EwRZoeLKtaKBntlGexSDZC2
NKVr3gJjlran52Tw6Oh0ELgvTxEPHLeM6jWnfTl3gjUZHN4jOXUUYuTp2ECim+JQLJmWKhPTZJde
2jXlhTi86d9ecbW5iA7N09LGPd8kuXJQ2F3t/e7BHWI9oGJGBC2HidvBLd/en/VYfcAsP/Cwve1A
CwZyq0yr59F9daJINaLI0rpVxg6+BV0C12mAhf7ls7lGCc4HdIwjhpdpc/fvwTs1pLox9eN7bLGu
7VZsqaHAHPqq4I04/LTwDRcqcKt2xJ87j5OZYDUbiytCpOvxae+SVXEQhY1qwNsaNBTBLegTf6c6
P+DHVsrwK/j4eCo1TNHwLfRPsVhLPz3NYRIo2BnHZEKXGo8z4ENRetvCPBqgXn1Mw9fp0KR6xiWy
M8LvlUc44+Db5NomSP0MDUwSfouvrZgZ5tvCxjXr4ZurK/O1pLXIwxWIx8K0xgp+jzIOAkmVIJ+x
z/oGF+1DprRT0dVxC24zkeRhpsPs9ZgczI06ee5x+7GPfXjR9PP3RPNOb68K+i+7DvRkC89qsZXv
rx42gACrVb8fCFetLv4Qcpkiw1ZPqCtDZ5aZENNN5bP8Gj+L4yPyS05T4XHUPjEWpEx4vYqeweoN
+0c5Qx3ONpV/wmbK8pQQPb4cCY7LYubCI1ep3xTX0yt3aiNrOyYBcBj3zyqPBi2TvShnoHjhJjut
75NUXuQ84jY7O1C8STyIxwdlGOIsz3iLBzlgnZfZWsh5+cBkJM0jk3IIMyONLOK/Q7E+4+4L61Iv
RXc7IPSKZWNF7TYMt4hXAXPBPNlD//CX4CEGqwrL2Lu0Kitt/RS8HytJlcHbj6ykiDQJyY+jnuUY
r9eAhPewPINUmdJtb9oQfiLXvIa6HAAiOzqVJssGK0ldxzi/ejxPl8b3Q7FSEhB2S6lC4GtmWipI
PTYqCyhpq4jTIEOyMN2oIJFUMfYjPEArmnwGrLp1xn6dX6vImAIgtLZr6WGmlU8JO7H3i0qNF0bY
IFJZC71b5aE41Lh1R6N7RuSUWvGtkHabu6oGrqjcm2X/vXbVutEiYa+LIDnzK35+gIFY3MROgo1o
e+CIC3MfQBA4o7/YPAoMCf/eiTKLTQUE+FZiL6uXE+/KNfjZXisaNPPAlfTHbKY2zLBSSr4Tngr0
XQJAmTQrEHkH+k8myNEAXodi1GABbLAsTPdrTeyEE7LACC8laaNoME1pkE9eyYedka/5AOQYTsZ4
onJjbmNYMg4gg2n47R2WM6EFHYPoTEF9soWkwn2/gMLJJbnbwcROA1y5GhqVLZmQ3P9EBMHowZxO
AH1QWBQYbNEEcF7CgDHH3OgqkpKzGWSHz+Moc7MHmdDhEHcPPPKafUX1ijPT+W1euM4+wIh1agIF
dt5ciw+odXofj7IDN9xAenWO2Rm2oaJCRUPJgcW1M5/D1TFCdAaAvycaH1gpddlsd+mCwHjJxLiO
WIR7h75g18Ii9AaEEMyPM6orTkT9G3h49UrFivfXGRgxrdYHK+y+YW4tgzbDXTYWBitGAot6urCC
Q4jKHWMs7hlMjBgl1RA4uvMuiAKbsAJ8mrQuF0N2ewsEanDpxi7If/FwyTCsAgvXlhj5ICNG7uaa
8Qkt7w2eYFumzjjtskNPJnoS4CXRO/6MwM7qwMFLX957yyko256onhGPT/KLYr9PrCqv00Q4kETG
KKfmXqTsBM56i4bi+spy8ytAvS8Md4OCP3zzAV7vHtk20du4k3WjluU6+deAxT6SNv+kvRg7+aL/
6A5BvMi5CWThJ9lNb0S6S9JlITv/dYgMCDuIfDE+V0OPQivfEssXfEP03NQLqCaomYAZ9UZ2xXgO
CaQBEwPvhp6Xih9TkyPx24BPvkR5v6EA5CcKNft6tWN7mv6vT5lIapugRLyHFqtiwM9AWpQuB7Md
ZA6PzNc+9GFjW5chg4JyQ9oAd+/2slKNSb4gEYcgCWIiwfi1Kq24BCXfKk2xmcoGynJrqPOJobpT
4Hp1Wxa+hpiru+uF3k8n29KKzz+vlasEBSHStWpCXZVc5dPlZGHIUUVEmJy6J8SbIMWTpPbxyVkA
DoGTPcf6Eab8f/2Al6fnnRcOVtDm17L2n8qEFP1qJHpfT8Z7TVEkdsrzYiI6yWsQFwHtrcvVjbzd
0WNffC4mUq/ewGILKyJYP7YG5q+XTRe8su+8x9cq9ouMKM8dBmwIS6UYUTMdy3/V7ZKRJg/2SDOI
5/HZJgJhsjLRuKht4NFoHuaH7we//ldUFc+UbRzt2cLFYqGSXFIiMylDi+3aK962euqg5RfBBhG1
Ed97QaNZjR8EI0MPnqexHr9bD493FgiyCRVCovYTMAh691O108N6kuId0yb6yQs1fF4G8fg5QEBB
hJigOzi7T5n+GfrMluzpytClrJglPsYycQXr1dsLFD4Hx4jh6TOw8Dk/SLz7jaIMDTcShBJ7wZNw
1C/la0mNJsVWpJJJl1XIW5Xw0+v452GufPIyrr49zOm+yzKASlJTl4YpMcLDYWC3/55KovX3MTUo
4y4Yfa+TbHiZW8kOvP+3fhXJ+J/GNbEsPpAg/Ga+yWDWFyWgEI0ZtA9JP1cpca317eRii9nF4fv2
veLUeRV3+uyS+MsyAoeOQUhuQ7caFsKeP+ByDJdRLaZP/CaEjFlo16bi8zywQAHIP3MMStJgPg7Y
dcSqLdySkGDaaxgmlIFEH55HI7F0JosoqeZI+JTpxZ2KswYMGdhdzLP7wrGPWNVBYYRQoNim2q1Y
xuKWoFezfdgJi9hexjmjqsDQVgk5BtBKppRoljxBXE1fS4MxbsRwBs0AHYF0xeesg+VT0zG2HnMQ
hPKxPLv3+Ug9Xu6CxCI1I45MZPLmeMqwyIt+OjexQkAKq8x5R/yJfBwUG9wYLHReuE4mbNBBrZHj
401pswdWbahdGM5OGMe9kFG4pmyCn0lJWB2BTJPK1hFAZXbP1JVSuuQw+o21kayKikRbNOsXl6ew
evkhhPDEUCp3n7KeAKK0tP+CPav2LPllD/1ti5n5qrB5RrnXAGtjDn3DRLVk5xXPcf00cmnlumyR
ot8Pbl5JJE5iVxkSEt7heRimZQ7ULTqZnWWHSHvYFjaSGWiJsoiatF9WKrq1iJVQf5W1QuAUD8S5
yblPzgcp2JHk666txhExYGEd6l/gTtJ86XUFqf355OnXlr/4US2cCl6L0Jkw2TekmmBlA/tlNxuE
ZkehNvATw71/D7K/SE00f11EYxp0Ky0kXgZWteUp9PiKfOZH1J9sQaQE6WsLZaA8rXrcfWETShKQ
eH4UHCtWlvnrqsv3bC6Sg51bFK8ETD5YFhXXmGy6iFoB7Y669LzUoWNQrJNErcz+95NBSnpQHnak
iFa1Of8PvqDVy42yn+U+d6iUFS2lCXgcXDKQulO5pCRP7/KLzbgS/lyZQ492n4Ch74pCrrh5br07
Z+nwz0VmSEmGWIxVqHZCo9xQb2bH1GDDSaINQlsAcDfvlyehyzHJQVQRusPIelEPVDPWpRtBxd2d
CE1zZZBjflcKq5p5NWtABxo934K7aoGfP8c9jUOrM7r3DL+CYVhKIRWA1KpPssLSnM1hrDOEd8aw
cwHPQ9XsK7s7wqcDtkSu0rBL5FSIyiv1qw+eleFNNx3jbuzdyGuj2yZc5w7+jJQcN5pDAorj+E9m
QDM7+Am6OdUcwbgeXFAcCqCKme0/0SJVhaHe152jz9qNCQL1a+Lv2vbDFsp1nPjDjXkyQv/AQEzY
hII72ToA9bS9HqE16rUHHtku+5dKnBEchnF2bYEQzf75BColPZGBXqhikrhssLthkxdy8fDpYJYv
jKXPV61pj1j0kRQEHnD5cYJjFCzAoMSdeL+0DQLypxgItStyI3rwMm3GSX2GXjZGJfUrs9XZM9kv
4fnd/cdHrcoXqSqAneDa/+T4tTUGmCRH8fE+t+hjtluxn/rwikFJr9Jlzztq+WzbsZZm3UxFsgJG
N5bVquChg3EzcoVHUulJgiwrXALE+Yebaj/+BVmw53CXsrsvjceHpjDY/JESDTl2rnX7WBmslBNo
pgb5R+HYUm9vfW2bI9sIaY0KbgC2sSq+pHBdlRtgx7L10zEoeuP45r7nuNvt3FOtEPm1xw+JUOxV
zhxyqhK2Rent5RdfrybHwRk8A7P9X/8FQp3LaLvRW3+rJGUmb5Mt8v12Hp8sSbIOYqwnGNkCB1Jg
PVdR0XzP3UfnOEzxb/dKas7vzZpASL1CSJbhSW5FaSqvkFkNkOYfQhwz/DWPf6UmptO1q4EkEfIZ
UumiukViLqr7b7AdlaT+cF9iVIxRFB+1/BJjcBpgKbnzb7UbGEgv8/QbVayAVSZ1fkiSTjW8sw+0
VYZ4cdN+tYpN5pCczLvKhp/UMZvxt6m5ujLEZrnHtjwcXEGX3wb4JhJ2+KuP0narECPcU3NkRMRe
7YCWTn2GVlBaP358AtkuMRKlpj5AlgS36aqYtZJPF4inOyZxcadXGYs3JdsEvYR5PSHWszWeOVIm
Ss9uEIccgJFFd8OkXRLm7x7F/E+OMIBTUVZ05332oeGwXt65xzYldVPJyWaHitvTAcw83vFegyW1
zDRkWcJIwYjhLaGx5RSt2b70Et77OGoMcPrbgHnUPXmDsQvJFisGZmwvCq8/Oua8I2hndq1M+QA6
kD/LL0h9HHUD7UDHw3YAp96p4usDk9yIZRPwJ/csLNgzfJoPHQLDtqEqRNBMJRNFK8dLdlomusgx
s9L6sUvzgeDkCIcohury2r50YwRkks8vYSYBxiiVATQyZL4V2Gd+qzGDe7VUiM7cDPJ4nYVhPQzs
Ys78mSoZNDDlQdp4at7ZT101gicdtcIbYIwlOgYahE2btzQMSjTaiccN3RK9ELTk2XaiyiJO9H1l
bEcdQGXeeF2GTs11aNDmTSGtIMJZ6wlpT/ru9wSWGHzQ5P6ARzuOd4qNL/H84JLOfxU0rwcFtfBX
xYaxnkCI6MZ3NBFLnrPHk1h/Jheoh1V94Mn9DPZiK5qzUl2CZbm1jE/6GF/oFnflTwBka2lxEzLp
qIFx6OrjWbYB7K2h7pkvnFee0640AEQ51qAaJdcPOztI11H3eala9aNybE2pEGvnszoWdHh4mLG5
kR3po6CeF8GzVKStVtksCf5B4MYHpm03oEjdCEZGMqRXrDscxNEvX1FY7ulyHRGmO0nQuGdCz5da
WMSRob5Fs4fISqj3J2VRRLh/mEaNws7AQ8Nhd1qGUR5Xki7+jMYNF4xQ38QfTBT35+XYS9yK/K/e
iwoiHIll/Zft6NhnGyWrdxDsJX6nl0t/bJXVLhRmU9l8zD5oHu3bb5/PbEPadg+U2k0NFw+jIoWt
XpDAC7P7JwWLjEkppa3JZM33qUQvlFrOcWeHLWdpjO6qPxc4r8FyfnzamUdPeveAcQXrUkZqa9sG
pL/79Tg5ufiirSqoFwrtqcBV1cHR9fIIKY+Z2rZm2YaZakLo/sr+yRy9CDswxnTF4oVD5YSl+c7Z
iaTweGqb6CcVWPFHO2yTSgMsKSTiDC1ITWMVEnrA1eha0EpnG5xdI4pDI/Rt/lhmB58mbTAKnkEH
gmAxOiDkUAGjnSLkY7tzj4GrsOLwlOQk1rCNk4DqKrVtn8Zu4a8JIKXm6Q9xMLhvlvEGUxOyJk5w
saHPT8FgEGIaEMnYCYU92d1BWY+ruQogCe/Qdq4zDAyaM5l+rozFsqMTXXd2RgF10rl4vaGK7Ih3
54ca0hwi2jHyFh35vtx9zrVY7y3bmNGMXzab7QL0fwOaI4VNMuDJKmzy0IGYqck5z6yVYcri2P5q
/oCtwr75p+mZP1dTBYnGoxJBTKY73bgNwxxoDapcYCDtu64ZePrfhOjXLvezW2hvR379FYV2Sf+m
HcMd8WpFTQKctoU70hOKEBHsoMsL8UCgP7xO68d8qiQleh0jSZFiDsMzJQHbk14CLAMkAdtHQhrH
losuky3KblWdBI7v+YH6lWAvd/vR7heclJQxqtUJbn3l4NcCkRMY3jWYISZk2+NEI6crkP2MHvMd
3nkoJau3RLKj3iVNDe1jZh8GRgHqLE37zsKn7S5bkr9RuAF4oeey8GPM/PO3Gfud3NDgFTRymqUX
KCAqVulhSUnQkMe2wUb9rqppGC8c7FnssUge6JG06WHlHNbLZlmbs9/UrlwrEL/56Au7S2BmDnHx
9rs/Mrt8hl2yWnsHb+Pvljk7DUMaPsctwkgpp4qWmySniEf5/7KaQCV0aGfMyzC3ooPLcPrDqcG2
4S0D4yBpcdOZb4flPp3NfFbpFtXRsPHH8Xx1NMxXt0DSv6kP8f58SthbhnU5HkWT2QL44XQ9jIBj
J0VtX1eAfzSpb5gAuc6vXBM3UqB1jZ6+mxwuomrxw8vlenw+kkoXQRO+Rp4crTqM1x1C/ILmCA1R
mMWIZXGg519i2ch0IhtVONHWbOKao3ew2kncenn7vu/Qj0Viv2XtwrY4t4lFAXo8g7fX0jqMdFaS
mCe2LnmyLWSFjKkG+BlrjxRDcBUx3d6dSOT3DTyPyVGEJwiaKZGuby9p5c3oPyPn5LbVrKmh5/il
s8g13103Emcp+4ELM4coDSa1nIu1ViqUJKASJKCUczgkg4TGxikt4ivWSUmb+hLEJB4XGdMcoblS
XKEsJsR9E2nDSIwkMVGcrmu9PoQQ8AwfTmNvBN+Ja5L/t+JQ1HPveiSBqdcqH4fXfgWBYB94hplB
ekw/HsxGzUbDqLRAg5pPG4GjxiOiTCX/iqrLEHQcWb8+vItpQPCpm3uVSsAf4UxTI3ithGxsehgY
2qMeWOI9qd/jpydxy5pBeqtVhOr0WvEjrCvHfUG2HxhKmn8Mzr2hgGyqU1xCJAUbrvwkDMwU/BkQ
ZIBkJwcHwzHLGd+To91G6LJfP7hkpOydu08zDaHfNcoO+0xbLE5eRX4e/d1na37zVDQyZ4b0cwlA
lkLdXgsaxoH0izRX+BuYYsDqapwwzQ3iNaZ5Mv/CcMZFP5nggvvBUDNZR4ceCFvEjuCZg0CI0S6c
HmXZglahAGmgPEGCYYczQnkZx2Ib3diwdclzyfZibqAYU2cefoFpovaVQEynVAWWYnFy7tR/kUas
V/iDRRLy2g+O6gYH5ZFlI/aXtPlHCGIFZvAs0/LONblkQ4DKPSNKsC/dsRXnca+ZR536k3sUEwZO
SzSA+Av7WXoslRRgcqed1pCOh+q96IFpJSVkYybJL9IwBAN77OXeynkSsP7tKJeLYCGB6NyPhz78
jQnaMqauKMV+4E3AxDOqpDk1P2ISSXOfY611gQDSGlEcQOsncZtelSTo7hJLclDh2BM2s6IT+mMo
miyLEC4geFU0NFzaA3rPfBnByiG/OQa2Rox++0605/H1DQk6XT1ytlHwhul9WbJC1yRdEBoPHu2K
vyJShs3CHWS7h0anYxye/Uiprm0qrUTiwt+SDcfkcOhU/EUWHiKIbKKOJQFknSiAGMj1QbC5eCec
QdEQZ2aU12b/FZqzQiywwSQvoymu7DkdejMkUIxq5odQC+5wIeQGjV/mbE7+zLgtnckBauXHV9RA
C/2qJkw1MskCJCQ5TOFiirZ2MzT35UnMIpZcvRzl2dBavdRkhU5bOSY/eZQugmey2UvO5Zed8/kU
snJeTXgNMLTxGvNVE4Ap42VRjCV0vP+HJJf4kgjKviCwng89A3JKV1QTvtbGg9VuCWiUHFKLft0t
F9NSjFDKQlEUwEDLS43JzTUYtDx1IEK+xKZZ6jlKAGZG13v+pfuk+TKawIO9wxsFC6dy5A+fKbU0
SawnZGHWwaoDZ5dYcJ3evbZjpwIiaM0dRyXPBb3wfspo6QsFgg33Cb4Be38Bvo8PiGM4TL+llzos
GnN+6LUmOdhTNd0G+tUKpIT6u8SqB2//9ltvzkpjJwNiR2JmkpSVVG1YJoesVBl2lGyFRLHuQTiV
iBouZTRq3Hw/h8qZNdfQMN8eIxafDxTCP0GxkHU1zxuTKKKRZ703L8Wpm2Ne2Rwzsa9VtsfeEqYJ
IXGaVgw2on5I8mJoVOFLKYbnF6Q60h1qzL2A6wbripvqZfrHtW1X6Bwq5Hr14uK45z55B4I1uSv2
0Zz7tLkIJT6Euc5SD3Jek9p1JvdFhj7jPXnnGpjkjJAEFu2Ico2XP3FcUNBrlH7VG0pE5dR6dSRt
fkfViWLmKG8mWfYHEnHrBnMJ/MsEQTXyimdM3f5JGPpiaoh31/BJ+avulid59UYX0OIWRnaAq4Or
fOra7qVavSf53C4DjZx3KmSRQIyBNTsleV3D2IXe+E1qVHRiSi0P1Q5El0pDIKb/7IVmRHAeogtw
lzopp85Gbi0o0PBQoOO0kzfuat8qDgS4R3dlzG4XDn1R9zNerN9J+E/NLurqFtWMNW0XUSgD//8z
LBvKiItrYO0AGzKD6uU4z3n3R6C3FB+50LuDhaSwAzqICQCmTF7EDgXbsDCecwptvWwBgSMjIcaS
o1BDHcIoysVNncWr3XMxCp5SCPpg/Qw1S3bnd2OQU6JoadNebxKhLuwpZOg1TNLhjvoZwE2sOKg6
PJ5ueKYEZYS8XafRW0Gx1gbbo3jum0QDyyalWS4leUiirVSNXXMkmQfI9bZXKUfCG9wKAbQTRsfU
/uFcQX7C1GPOWnBm8ScNDy1ko3mE6YeOeBqm2oKyo1n2+RkXkWA1Rgw5WGwYAAB9RqwmwnmlxkiS
6sLqwc6+bGlob9Vl4j8yHNXWJlyBsW6YuFx+Ahpqx/3Jtibg30Dgcm3vdNsaOiekX8qajmpg+eJI
N4b4W7Or0AaKh3uYLxHFO3MwRppLoTXZLcne1HuMfSk9XYYMrNyh0yG8mW4f2hdNhRULkfrGrm5N
dlcjmhgjkTtJGKqoxKoGrBXkUnlQgvqqXsM3BXLEh/xZjRqfZ5wRkpE4cEWDytR8a73S8R37tsF/
xTju/PDQKDwG0wcJLp0kZG5VeBTJmzjPrhzwTBI+uKKwLh/PKgUMkNKwOfPI37qbbSk5SjeNJ6Sd
DZSVamJSMKD7+y0V945pLaA665apl6RylV492gFv3YjkO6r99BxKJFt6eibpg//JX/DzJVwo3fQ+
Ek0GvLuhG5UGNrT2A/CnJNn3T+l1jlPW4IL6z2XYCHuqZeEcQ5kUooDFStan2M9zBbULv+sXEp9u
A1t8o7u4AEsVnCfzl+XGYPc5UmIPDwGpsO/GtLfZpIOEvcnJpjXqwgLCM+VaBlJFMp7snIAeHgxu
/4yuD0reG1fMRyEpytkheP2UgTNeb0MGk8+g4lec6ZQqNLKN5ci4MB+d5VL5z276l+G8mUXpUbXL
dH/7IR8GwrqNK9pZYFcebBiGNYgKawOZHmie7qOKX4Bxxphc+RsSamERQ+bKZbYGWqaMoKqa0ysL
jRWldLJXitJ8PErE0bJS/tuR80W5r3Ot8CvJCdw4DvEBhMHP7C079BqDJaredTc91QJFIPd/WUza
lwhcArA3PjbXfQFoApHk4WFYRP0NLXwQY6ZDgA6PqaG84r1uOCvNaeNrwbBb+VYxiMRH8vmY/Mq9
dYt1kteb1p+d82w8PtVKvblGna3vlBKkXxCo8P13EanxJOTthdHDtVSngY2E5MadQgFvFw/WSD5w
/A/RkRMaZ0Ng79r85BiEnZkYyGIfeLRKXqaBbP7UtzngO/daBVpuwjyeKtK3vI+3drOXwS1B4nNY
Qv1knKZUIu9fmzsAQcPkyI9yBsYcNjDceoaFXNreXEUzBa1TrtAAV2wYrvT+zwISxrmm5Y40N69d
rm6BB815DluEqwM4Z14qWyhN1xysU0Q8GpbbV0FxGL+aeHKArh+fooWkTBY6+9xS68aE5IXKvsmZ
S07qzXQSSbpTC1t3sbjMN11Lv6i5tPkqk6UkE5X0+bWhXIK16ZP8oeIswewruspKhjt3OxB2gFjA
wB3sDmC5Xx404VImBh117T6PUxQlDCCe7FirT6PoaC01rT1fmbqwOfd0Pbzf+RrPFKTD+jjH9eQH
JsskD6s6OJ7pmH6clYmJQix02kFjzFPVzOq5lLk2o2lihMU1WU1NHuU1Ny8+6uBmRD6FqDZynX4a
h3R/FOu6MEF4ScPd7KmiLUjUme+Nz/PQk5XgLST+n1tsoEy6m1F2RGfiHKkgxNLmqvdtw01ydpnW
NrJFPbbow69h7zpc8iTmeWF/clDxt9mnouO8NT9sab2nc842NNEcdqzxM2b5EPjPpJ1YXFXfKBNF
/6bHu12t//QqMzvGKnrpx4D+SMKV8tNZZc1kng4iunf36HGOgC7UchsmsfEgPx0hj0l8I+KpyGy6
+Bg3UgV7eu++XqO2sXsoz6KwKPFw61MBEpUxMYG765TiGwQTzkM8c/e89QlVLrRjRQDDNNoSly0g
SWqVD5NyksSRNoSFnEnb5UWJUnk+l30lhJy1XzTkdeSbBtOYdirvBcPBmAfpMJ6kozmhY9asNrlo
kYQUoKhwMT4PILJsi0symf6AlMmerRFn1UOU6XVY9QirESv//vHMMliPgBTduJ4u1vyFrnUwD2Z+
VKb2LSGQzLYUM5vTgtQKR6e0yY0mXRS2dDu/rFCEnFCvcJNumq7QG/RFEgfKiZMCY5nauCx45mVD
OmiLh7/jiVFjS26sRMMY4OSmHfwGAXV+S+M/bdPCHUhVohcq29MdD/fAdF3kRTEGuVcGGWx2AKdf
SdnL+YIdNKyRLkR2R+595NT9AaZCQUqpXiBPwaTjhwyFJXsocHGLN9z+w1RoSz+eRJDc3Kzfn38e
f5Z1uqlD9zdn+QCaRCQi9FuGtrAA1TP4AMLbnTkSBINnkbz5vvZrlkO5kgryZq4C/R1VMVsvXaJm
uNqImJ1O17TWNeY0X39TJJjCcVIiLnjg/YYfCJDdHB4iwsRzIJZEqKu7OtS18F3vst2bJD+fA6Zu
q45IoB62ZH8oGMtAh8ahed7sHSM7uOqXw2hXA0zxOVMiVdcM83z9Jo0otu3HYhb6NQkEFaR/VQNb
6SWtNMtPLYUWo9Vuz+3NzEiUe0FervOJSxa4CeochY1URxO6/FpwfL6gAgsAUSnyzvVYjWRlzFVS
hJPCoLiCSGQ0gHykr07BBV2oPZhyPVl+lW0+9Dv2N9nqQOQiMa8BDxkLNMd2yCKYkF9yOUzETb7e
Dr0o7KXr1vcwFh4jTzAmV91miUqGbuVdHqsCh7BAYSWcdNamR6Kgw/Kyc7IHCTAEsdgmYRGONueA
eRs1vSZl4d9cmJGtov6B3YW2bd+b5JtIVkGlf9w7Sv/ImJziOvRJzHspvKgiZ8z18kdf66Es4+2b
x8YcZXNkYEItTaen4AeQ2x2jkuwmcGixycGIreE1EPd6kLPU4GD32tzDH+vgtvbLHzpoW/UiGH37
3ocMhscOGxmJRWugN1HzAt4Zky1Fm92ifrb3ECvZpDWOCW4LyS4Bo/rBUqBFWpoZHpqzSJL9Z1+d
aLB601q9d+xY0agN2CS5whZxATCqMGof4wXs7bQndydT5GiBdQFDBrMy0byENngsR8gypgWeiRb3
y3C/PWcC+VIoLkKFjiHce4wbOwImyBcmvF2tVakYOUtFsL+PFfEPslYGndoalgx+Ih05YastrbhP
Qkf30s8e2TXevv7EoTvZl/5Oy+YofigyiN3Bkk8ap2NqnjVQQTHBhPnX4SPZsh2b30xd1sQxfJ/V
37xmBGXq/z1nQrKn65ED7j7bhuMu1vDRZ9P70l7gobpfl9yG/U+4NMPxsBCVufiwDRwm8SFkxy2+
5NCNLNdSBkl51NIAJMQ63BZArbx1eTl1jIrf64NMJ1RjZT7EW2uF/CN8rLRlXVepfJM8K/LfKgwL
n+Zs3Xe7qg//i05xLlDmq8vZw+Kr1qW04iTlbavkD/JFdZgc+aB8Wc78GKesArj8XZ783Uxo8Q1C
d2CT5jxGiBJKPrws57hIt/Qw2zrBofvYePYdgZ1tiaqetdp9pRtzzs6N6VkBzZAGogMcYRhvTt9x
KcGt7kTq9ieSD/8SBbxbjxjk5TqZGuuX73rSO5QSpyqn38w2gEiPJpKfyCapIxRSvv24Ze4bJwvI
v9EaHJmDToKVbjeE3o/lUTwRTqgxOHRfH/iQA1oEfH+sMfJi8DZib6vFGZzAuMwTH5HwqOXBmQNe
kLWWvIMm8NLES7Wb2rMDbw4gfcUVQOHUjwplctLhcL/MY+5EFPnYvF0p5DvPvsDMP/m0SLblloAT
aJh2iJkXLYFi5rOhxeB6GZatQbF8BaZYJ8kbl2O0KtVSTnqSpaU59kghyB+hCD5irHvOPN/6K1ZC
hbx2txQVnZKUvscl0k/jgg7FuPbz6yZUpUEc73aZLUauzZ4LzxyolyArPXk6h7DNvVDQNx0kdoIT
aR3vAvWa8C8URx9DnW16JhN1jJkTy878exQ45tC+68xoAOEvLIVuFL7nrFjJRnd2ptH0EWmtKiqS
H9XV+yw4OtqedFeBsncE9yCL1Wn0o53GM8JItuxlHHDh4N0i+pbZ/wN1u7bc/JUtPoxFA6V8DA/+
LXO3cLmYbhPDTsYh/ur9iXrR/6kv3oqqcSOT7U6g1awSLNEyrYPzzLb/TjoXQPUGSpXGOba5coMQ
Dw5M/5IfTej7G41xyLnpXnFqXq066Zk1V8zdVwWsmXrq9IP9UfiJGc8RDUPwox0lGBkSkMEah/tU
8oDZu4RdHX/m9HuxKEJrg9uJpFy55Hzg8942etRlFEoDrKkBbyjOg0nD5YW4P5HzXRomwkdAZMFM
FYuvs1/J3gYty3QuzVaCwZoDKkApVQIMvtG/yrSbyWR5XZcgYYDpvmNGVy8O1JoDD1UHgWg/mH5c
WC6cQsiN/eqYLwWYqu+LWB3oNv4AMRWovI6vz1MpIoniTc0jb3JLyCJPufe/ixSgDniZlfxloEFt
+ioW30EpwC8byR3dcnYE0ct6ttozmv/JokqqYBqp6QcOmQYYwoR0UicO9+A54q0qcu2A3JLSojEE
KjF5Ofu0z/fSpPPEKwbCdCJh5M4+5tb+HvM7J3z/8K0yn8Qm36OWoKdFqY134qJKHopJCT4Fh7Ca
Ahv314LkOMH2mcCTZe3biYHsldDFldKI94+7NXgw3AhSfJhCYwz0DO+tj8HJ29t9dMNJ3kke8EmE
l1YVdn2Pz1xrmJ1tTVaLtzCVL7P/YaGtirfVZz1cSi9kQYyJhymP9wySX9OFp0kDbHLFpzF68mY9
x7RGF+Q2ye/PpRhcONxe2yqWlZDxV7ytRzfRrAXiVwiZNP72ldIm139Va/N+st63lX6Urd6S9zk5
fL6OTpN3TbKYkubUiNpQxB4pn20vIcLyWGV7TnaHq+i7ase0+wQKAJEFw7iiLaopfF0zI4j4gYs4
/JZ2L14sCAruZstx4LRds82EKtwELcaTEd+cqv2iOZj0D5fhVbYueW5g4GQd0Ertp21uJQSibQry
sjjGNkHNjqKAeALfR68NdQH+FI/UuqX6XkkrW2FbV0Ako9oSU/P7z+jvAcnDIT6fv9z6P7zOAC+o
MqJpQ57V8hSOQEndjfRVO+jnFq5hfN2vgVbkLiFHRHUYUgR4bOu2VeGLPjzqMV9Jll0bHz4Zn2mD
2VzPeyu4MrQm3AiGjKa5gscg0y7AA4EPxS5ZDEwxHCNCerbICA9deQ9CHe46XSotn173KlSNcAZK
BiJfWscQp0/8JU38Hprxm5Y1fAlQkl6kpIoRw919f9UCyXdyuaOkPzpqTWPPQdJp3TJDOIn05nn8
S47PmLJV3sZX5UXvDZXS79jIJW6UxPCsoVjmqJHYgISzqSSQu/R15iQI9c+8ud6r5FIVnX1N/ymv
NI0wzQAEMwMnm1+60k7Ddm2qzKAQVO80eAOXZNFZrbGj4JLMNoANdoKFfyTHh3vfbpJjROSADw/z
U16tJV03HHAoiT472//jvnyJDByUF1qfUZTHs85rX0bP5975BG1TeOX/FNMOk8ieKG2M0dcosUQ7
eG6ba/dKmcWzP9drtRmMqenFnVPQAdCc7tNdD5tS7vOtKnXmNAuSvc7Dell430Tq1IzmfpcacU5s
IthrW1mcIc6BxOmw/KmDq1nUOAbR+hURH01ITUTqb4pH01POJz1nzbEdbeFgdbimErAfsce8xwVT
RcqiQkiTTbA+uheD1nknrwJ886suo48JVJWKYYJYSdxTS7Ibj08dzFQtWIp6QNKZRw64JRkHDdZk
VHiDmswTfK8WNtGRl/Cj/fbLqlNohqoti4qSutvnKTgBLBXPJ2IOXnL7XnrTRQsqixr5rXJphxd6
r+OcVczCVI73w2B+eG1+xm3avX8qltNISwpDvNxwjYr0JlA/wTZBhvBoomo8qZMbE9j23R4k41LP
XF5od99Yf/LG0oa16OjesnKqAiQiaKQ2tIY0QIl2gCZA2HwmKgqP5YoFy++DrJ+7lI3hEmhpWwqG
4BJXFZYwzNHv38oHqw9ZYgLU1XXQw019ByMbmGU2QKFojhYCk2GlL6A+sm6LRhdbJzZsbcw1UDwc
NAJT7LHizuu3RNi3IcfCqq1RjVeoqbHJKugTvuAgWBOlaoUhHIJ2ALNfo++txClPfML+MT/kgyCj
wT98R+9JZ0WbSy/3+ezrpExvYzBn6a9rz4fe4QyaP6YNOQqKPi99xE0nL66KVnuUvgLss+xEBGmI
axlPRBuaNv5MflZ5u8Xe8pu6gQbJU5YZWrB3zlWkzxed9rNWaetOSzGy7m0P0N4S2q6NgoetuzqS
rDqCpCpT7bGBwDq3M7yox5SYCl2/KVoeFcch499I4RZIqRDwosg7eC5t2cgj4AYXMTZulhMpTwvy
CVf0xDRDRLCmVDGbIH7Kzi7ZbrBPlQOyBENgPN5t0ZNc+I4tcMeeKlPuMccvpjZIXKgrlfVRyiQe
nx1ta5lnw49KiipnTVwEmVELY0uWQRx/pR9MHNdQdFJ4Bq8qRXrCZ2EwADFh89+wd2RYgl9qNLfl
8BLOMAUnJNfkG7/uVbX+L3qF7MB3LJ4Nf2emRBmQ+oVygQOR91UmLos97gRU+9eEYYdCnvkklZVt
s/5s02FxNSZ7Gl6phr9x4fGUKsXafJ2VxOMS+bt2QNf8aTt4MtqTtTAZIVol+BDqiCQWHbvPr4nH
LSIcdpo8l056jLrnKp2EIg2Zh9dPnzwm/PJmxg37JzUjGQzOGemyOWXSwWvy6hImmAtHjXZNHigh
dz3h5dSXD2Bsiw2xPpSlSU1qW3efH29YJa0tqaV1Bh65McQQy3BpXvdCZpZ5+ZiMdu3BgfCMyKxn
MCzi4GOOSjbA3d5LPed8i6b1YDjTDmw734M5mbSCfwjJ/NczAfIsUbruqJZsE/IyxPrchidLhi0m
7BVzprMitZpYNTLs/a+9cj8KElRiW+bH97iih6YGORNYmsfCvnE9ld4wjQACV97Bfnu08qqztYUw
jTxvutIzicqcTNMjM4uZrikw27FW41UyodFNaTViJuMmdUMED7BUVSTx+AKhamZLeH0yp4z+JMEi
zPbhrbqqEvZKxbz+WGTayKSQ4K11bBBwnlB0FHJabVe+oHVAEDe71AQwLQGKIIOhytDKtKe2Ajb0
TT/QrK+7y9zlUUbnW86IH4R+nNmu5nufoOSU9RPNqGp8drhI3sk9+4pdItdICVGkLrAD53P7hcvI
W4IR0UEubrqJiWUEwGDurXcFCda9g15hrcno0QutKUP1c7DpcstPiJ+4mkstDtXpGMhxxfjVLWNf
EgxO7n0+zOkZ7JqXhuPnlCkNNclAMRd6t66GycCsvc5zlomSt5z5c4dECzwCli3814/h5rhMLfcU
Ih42b1Vq//nQz/dU2mp0enVbToQBZm+LYmH5GxKynN2KjkLK3o2UN0WeMf4hAFpnK1j5S503dnGn
tboz6qRxynUvkNZQFlVSi3iZnpT9Lg/a73rVKKhSniPUMRrQ8SaHw5k2LIfT67iVLyIQU15EoRnN
2YJwKAI2+7AxfKyae6QMhKAC1gqgzfz0TGAfa4aWpjUAyosTQxun5K4O/69GYNpuv0Koykm17rFM
/B7PhiuxKvZTOKjkx5DF3DveqVzIOFdknUCaupbHrkNVFv6yVTRhsAyYBrpkGpAODTJ0ymvVyI57
Fp6aEvMw+IjCEgphaFJV79Zte83BlCvhVDs78ByjndySILMa1gNnMXTItsIwAJKT9xkdj5upyUAS
PzVGd2YuWJMj1u+13DG084BWhGfnRldj8bzd0jvquWLZVVjP3h4GrEPFwLORzp7zEHBFU3Kv09qL
fwkqhUVxVXEtFXEHRC092hxMan1YnUuLpf03msGoiVTQB4GvOwl3FS6x1qWjGYXtVXIZBiiGlcst
G/Z2W8Si/7h6bf2MY7DeNQi+HoAs1n44YCW8Wj7q1TjMymrKXH1Th4wIbslnHcR71aIJvLLXBOp4
bogeOakqFEa2RHcMmvVMoGrsPeyNn6MGTgjS9CEijSYeZrTyPxfwRzyMY8vBd8gweZKIB1TMEz1x
B7sQlzd80uUulUrjdOX2kBxlsWxakKEkWc8oXDsTUuqHy0ZCOwR/SCCnjFTQorpDnaL7kb5uc80S
MJuLdF9hwhKCRY2uOBv59ET2dJ1aPnq3mpSG8l015LjyAqAnGSjCWZG8c3oXD81lrjxPZfznP7N+
p6hlFqktgB/H9A+iqiqjGsJLM9AcE17s90JjyLA6/xgk3BI8r8gGxFOmKmV1CYQcum4rOCO9MY0r
9BeAfsmqm6UuP8tp2tHAGzZlNdja4lK9V98K1ivyH8XcQdXImfftJ/obaEA9CCfp2Ie9Ld9+izjv
zyUayL4KWxMenhhacIAB/Z5F1VtCQHRd//hvpKBp+8id5tPs788hr4c0fEN8MGD/Kb8oqwxZiXza
Ykda6A8uaqKLPlAD4zT5JoCAhyc12YKqvlgrCcsovEOa+Ov1RyLwChheeyOnoFqF7VIQjWnv/xw8
7+A0OoKodS+jK8GCznLw2Kyi6+TtSNmmpQG/I5fLRiyUYLUlXaN6n0VUFjh5QcrGd3RovrejLEpZ
JiNXWkkuNoRdxQblX5XFWFbMdHk+MVrsB9gMmZps8krCNj2yY4v1ayIzN09N1ie8v8Uys9ekDph6
o+hoUjiVh+k/9VR8B/znHnJ3XtjRHlK3rHIklhxXkqsDd7zSrpM2QTV6bNQCc7DACX7OR118GTj3
/1bPhVE3umATJDU6k0RjNMji1kmRfccBi0J8yow2R9EiOeA9RK8VVt7vmAk5I99W/rUnuh/7aEDC
jlWvUyz0BLEfb4VlzCzLUw/hM18jGYWltnztzMiOtsj6Iy6MyryPoGwFpozJBUHZP2f4WVQeoyA5
Lb418VRSD2B75B77GHUvGpyY2/en5BG0p6ZF5u3kZLMabf+W1CGvtLKp97DB7ZIJcP6ZnVV+PxmP
yTMvUYX8EJw4gmBULALWYXqaB/2yGSKknL5WeHJeG3H3vHIXiQTOmLOyiTQH9ODEHCV6s/w3A5/h
MZQc+eoahcf59xcwd7SvfgChS49qVtRfWWkpMRdnoN/GDeqBpqJnz+WGZL8KE99OvcwOfFhsSgs2
1Ri1ypSr445lQsaPqIosie1S7IJWUJ6fk0pHObXJ1gcWv/yxDfmzx3t77yaZ9mq8f+XW4Q8sHya+
fmJOpamUNnrD9xIwCy5vvHmF7vi3ZsmltD02grINVmhTrbEYvfbk1dq0pd4pG7DMerVL1yrkOfOP
Pbi4m/OBQVOOtRXS7D3QQsc/ziVMZLyXbzgvOg4Cre15UKsRXHLIpfEiSI4uedf4zYWtShtxzF8i
RFAwG2q5T4/49MBPOTwemXyPncTde/zKhM8W7PwCzrQrgqBzCJj7M9b0ih753yXO+JcFQ7KG/+S+
dvgUm6MGOnPfwCPYzCZ6DBIUJGMmbAa5DQU8tcfC7/i777/G2OLvZVfBLa8vQWIoBbbZXG8g+wpM
VdJcQzYukXFjDDh6qJ5lrGgfiUOEKJWTpoFFUX886eaQnzWEN3+NhMvRohhtu9uqfemfJjUtRoIF
UBbeOJpGX3qX6ZL0A1YPzMS/jZEj3aZp/C5pvPEqbGSkBXLW+doow/NLDL4lIeB9s6NxOp5MlvPo
tOtI1lJDflgD+0/U3R89GLvv+TeT2RDqZPPSRkfgcbvSsE3ujhy6kOpkJYWJB78n35S9qtmIGCYn
JjbbKuKz/2mpNGUXFnwsQ5EL1YNSILfwEBBKxvQXTiqcLF3RojSFn4jNR0Ct9yL3elB9Eg7CJhGn
u7GjZmAkj4ZUS1+MgRTw6eUbFP21GprE2AIytm3RBAGYsiSIsxYRTCY92/vTt0R8ZTiLxHthLP3h
blQwUtVlkD5oVJCdfdUsjMED0bmQyxQZlRvjnqbOehF2MCU7MOYzhJWjKqVsQxSFiyZkXg7H7+nc
cEdDGUvStI+6+29hz5LfjwAQrn6gsZaXKDhcu/nCbtyI0pk1aYV6oiWKfaJqLalILHt0YUmDTJT4
K8yfML5cbD1ToufB85MWKo1URlkO/UlRKR3bR80LVOH5Xdjm7Dje7pNupJmzM8Dyr1avSI6/tKcy
TIXfZ0PrkEXPcDjpG5FFUTItPyYM38YwX4agN2/j3AlXD1p0DuSNODtgjYYGEm9/zbCajIa7KuNg
j0eQ/lOcaa2kNuKcRPHZsx7TrKwIfEgMLDCPfd/bi9dMSg3hEZ+wHZZnitEPxKRKIxt38TrDvC+r
8O2GtNqaHI3pvV1czHueC9mOHBVpfJxMXXceRMgRVxnDDc0Ynkko1R+Xz6qzxlhaEpm+QEONqeL0
K8wdnGHZQxaCRH+lgNCuAnIFvR1qihKv9qRHucSkT3uCtcwi6F9DHXHxnkm7FIJTAi36E9+GfnzR
R/UzjjzHkrYJcCmi/6haLPAMLzW2D2J7LIhAqmrT6ytnF0m7LDO3OseCL12zYYjQOoCytGytSq1t
2d7VqhAAp66tndt4zeCLnuxWmplqN4EyJReAXwuMwD0e1NnfkOv01/hNyCw/O7FegMbyUNSLjjPm
gg/9l0Hn3+wrsryQPNGlEB55nuHt01pnDsw87HkBhUGnkdvgHiO7+yIJQ5kQXFqvqdyh4mQphEow
mdnq/WmqsdsFc4zviT15FwylsekTGcB8gE2tZMCEPaOnr71mdRLQYxVbv1f6R/sa4avv/RyoR/AK
wYBp7dOKKwM9CO1m2aDITpg3vJfDyZkveLSu0NQT9Loq6c0vniclKVJr7a/LAyuttrosAxPTH3h6
DeTDWW56q/5dWOxqchrMcmEKeqLFirNtVyjrMT6jraQ36VyOyA3iK0FPrqWgNG2Bnv5E5hhXylno
xJroXORNYqBmOoQLgs0ruwMLC9EyBwrS/lLm4Ny9vi66Qeu2ZDZkzam7u+BZpdWo0j3Ot6bw4fx1
qeiqLKiOZXzZG3CZKd9qOA5jbnIIYhihfQmxtxYuRV21JN8xV+WGnp2GkpPg2ywy6pTq4ErAjr/W
rebQJ7eFuppoPk7tN5LD89JGdiIZtM+VdHI5OOX8coR/zkcCTemDMlYpw7txieHQWZxKTEmNvp/q
Fap/S2jt1OMohzdu3f1L4Ao996dDDD3TxJTa+AFpw5+v6m3PTBVX9l9Ic/krTHmHml524i4slbel
qsGF/lmtLo8bfCEovZvz32M0seAUOOUFypg6v7sdxtl0+z1b0NDM9jXz1h/o5DmCTRp29AKKBKdR
G+dmfef0EeaHL3FksSTkPPD+4ePQZb4f/ORPbmREQToVCIbnLkTpX/AlQ/YPsC7NPWmWiX42Ur4T
XTybvgbSeIxQY3jWZPLPiRSZFD3pJ3efH/jZykucAKdntBIoPfIyN+iRM4wzu37Ae0+ANIxTnGRD
8YbIK2mljWM8E5stvzOXNOR9RwbtzfF8O/E3keuQNqGutEIaDnj0INqdGgAuLACAyURJGaHTiJb6
AH403uyixa3y7OVltJMya532KUWouh24d8u2yA7XZ9r0IekhV+97AHGJ9AjBAlu8cdrU4/ywAR+P
cdn/CT7rcwzEdSUb/yueIDUo/R9YPt+NvmUq6SqI3g50dv1fJodolSUxCZd++vT0d0NoGWIheaN3
I45aMIHL8/oee9Wf0OTDj2I+hmd+Vkpz/gGieTQMbpABRuWYLVQhQdx+XSy5AnNrU8E4Kd1Fkj7A
36iPNzISZP62D98w61jwH8b16yxmraXtNakuwDeXmf0C1vKWCw4Qh1f3bUgkJz+oewiKFdCnkLth
I6MDUnM68TRJsMWv/WnR5FQEOptKU7clS3BfWpsHxYT3LEM/+oSHNd36I2Yi45fJHgVTq4HNoOoi
s64StQvQXAxfNxogbdMqbBc5K0UfirbA8mIuql5r+XBj0DIUIIWQHjB1jI1o4Y7XmJHSpTjwUCRL
7REfLdf5+c9J++jIjSFt1aEjHUlC0wfw98DpGo6j6llRFBNALqzKxJLU0rGf/Ao4O72D4uPsYJt/
lmO8zBEuTWseK9dFD+1Lbs4RLO2kYs0CCwKXu6zATGzzfq0z7hOAhtdO2SqWe3qDtUDPnQTtACc0
L8DcC4kO4IKQC04P7bOVc/DuvBTGe0ul1w9ZHy5Mw09YeddjREAKJsgLJBu1xpueyE5MOhAgy2pI
dHGzUZuDnVMZ6qIEbF7PUPkiRWYyGtBwpTCogUR+cH6b4J/Mzb7arMZc/xfmg0OB4BzRZYZqf+OK
mpNv8WDoQPqN6tLE/zS5FI561qUUpDsjq0SJiUaDjG8FCtvektoL6K0A9TNBypun6rElVvN92QcA
qnzKE1cwLO1be8Fm4FUzO6voPtl1oq28jNo9Bh0EWoAKk+qkkK7ZmEqLB82cK6msUNNHxSIUf/dJ
LvjzzMltHqkCpJDvxpM+u3wT6/y1qWniR1unAgnUf8id8VgCycscbL2QC5JZdwOZBsgsLv60E95K
hz7DXwQd0Nk3aXn90/p/5E42pXkxN7dl6hczludOPTsqdEsrx21MeMbA+5OYzvrW8utQ+Obo5wH1
eDxm827OvPPWM7Us0uO9Zejif+KPf/npahEFpiCRPr4/UomNjimsfm9/JF0xquUELxm2RN2xf2Un
TV2+NB0DuTWOOKPjsJuVF0St0qkVK20HGrzQmV29DO2PXgEXwgVVsos3PiDm2RZG8OFJ5GGwV3jv
fzyuncNO7OyibfkoIX6k6yPpjc7EgbfemZars1eP9kcZUOx4vLQRLpdwtaMJCo2/cDLAww31HQBF
ufJEZWH89Et9WQqdjg+WVfpL5rqJsKexoRO835WhurLFZgYRqHLSfQtoR9Hzp6GotNTXEUEDky13
t6SVjxRWEA++Ri4VnsUhdao/iWG1XszU5sfIr9Mt6r9gNMMOMuQz12CYgoWmVQwHNbpLStditvk9
YINvEGBgOx34u0G9xPOLYThtl38+tCJ4aSGiftKrKtlyr3HzSqn4tMFBQuQyrvjGH8jdy6+No8B1
SXATT4udzdpyiONxyRkOATAazsZd2NqZTyD3v8HFVO+bXHrOumHCYqvJHQWrxQ/vZ8BL//omD12y
mq0SNepKqYombvUQ9xkUTEMyR/vSM/XSe1CCca2tevXtpJUs2pY1Fyf/k2MXpyEy58R57+nmcMyO
co66KRBafdpDexnIFMBXh4p23Nnr6NgL02w2WUkS3Vwx4F8pYSQUbdrrSzqdjF5MR/xGj2BHVBYQ
SOjzM8emzCA/GjE/+n8LOX4ndyGe82kuZdkUuJt2fZsLeG9m1avLj7Q5K9NcPcocYu5TALDe1+5r
i+/0suDAOfJTS/iJKVgG0yWFYGUwfFJwLCHOqnEt6c67TRDha8pXGUXxR6sWKNcM9bYXbCjYrau/
8QUpBi1DotzdW4GR+eDE9i6FnZ071J0jpH2UTsgqh7IStPy9NKTZ29VvK8zGj56QuVmvYSbUqNVa
mI2JCHJw5J8bmfJGpCgxupaQFBgMuo00pAz/cHXZ5CbcDc8iSSF999UFMTcOTg/RIAaGcH4Tm3Ni
6lK0V74rjs//CB4Wy63ULoP2b7kCdZwm0VGdrSnmk9UM4ao197Ax6u1NBKWtrXux05fiS3E534nE
0RYg/zYJxUnccej9TAYFQQrs1pWQ9drahciKvZxX//2B6rq4evg1jIENFylOyoVUrd8y2z8pzQFw
9gPgburXhcGI8AsUNF3X7/QJs6jvix/tX+SsxMDN0+LvSuZ7T6+b/IegCgWyruyv1S58g1LVJP6j
rFOW0Mh5+HaURudcHweH8TBOxjyuK9CsmviWa96fhdIxIi2BnU+ZjCs7ahO3/nr/7Toftwq6oxbo
w1s5/pY8Et5KHQibg59gWNw31zPpHy8CQEZ+FlS8bOC+C2+bOfr7VJTlUpkLk5DgD73joB5kXZr2
BRBsnlS969WjxiMQt8msglA=
`protect end_protected
