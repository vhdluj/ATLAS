--////////////////////////////////////////////////////////////////////////////////
--//   ____  ____ 
--//  /   /\/   / 
--// /___/  \  /    Vendor: Xilinx 
--// \   \   \/     Version : 2.5
--//  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--//  /   /         Filename :hola_kin7_gtx_agc_loop_fsm.vhd
--// /___/   /\     
--// \   \  /  \ 
--//  \___\/\___\ 
--//
--//
--  Description :     This module performs TX reset and initialization.
--                     
--
--
-- Module hola_kin7_gtx_agc_loop_fsm
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


--*****************************************************************************


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity drp_wr_fsm is
port (
lock0,lock1,lock2,lock3,clk,reset,ready   : in std_logic;
di0                                       : in STD_LOGIC_VECTOR(15 downto 0);
holds                                     : out STD_LOGIC_VECTOR(3 downto 0);
DI                                        : out STD_LOGIC_VECTOR(15 downto 0);
Address                                   : out STD_LOGIC_VECTOR(8 downto 0);
state                                     : out STD_LOGIC_VECTOR(3 downto 0);
done                                      : out std_logic;
kill                                      : out std_logic;
rd_drp                                    : out std_logic;
wr_drp                                    : out std_logic
);
end drp_wr_fsm;

architecture drp_wr_fsm_beh of drp_wr_fsm is

signal store_di0     : std_logic_vector(15 downto 0) := (others => '0');

signal holds_reg     : std_logic_vector(3 downto 0) := (others => '0');
signal DI_reg        : std_logic_vector(15 downto 0) := (others => '0');
signal Address_reg   : std_logic_vector(8 downto 0) := (others => '0');
signal state_reg     : std_logic_vector(3 downto 0);
signal done_reg      : std_logic := '0';
signal kill_reg      : std_logic := '0';
signal rd_drp_reg    : std_logic := '0';
signal wr_drp_reg    : std_logic := '0';
signal not_kill      : std_logic := '1';

constant load_addr_agc     : std_logic_vector(3 downto 0) := "0001";
constant rd_drp_agc        : std_logic_vector(3 downto 0) := "0010";
constant wait_drprdy_agc   : std_logic_vector(3 downto 0) := "0011";
constant mod_drp_agc       : std_logic_vector(3 downto 0) := "0100";
constant load_drp_agc      : std_logic_vector(3 downto 0) := "0101";
constant pulse_wr_agc      : std_logic_vector(3 downto 0) := "0110";
constant wait_drp_dy_agc   : std_logic_vector(3 downto 0) := "0111";
constant lock_agc          : std_logic_vector(3 downto 0) := "1000";
constant endstate          : std_logic_vector(3 downto 0) := "1001";
constant resetstate        : std_logic_vector(3 downto 0) := "1010";

begin

holds      <= holds_reg;
DI         <= DI_reg;
Address    <= Address_reg;
state      <= state_reg;
done       <= done_reg;
kill       <= kill_reg;
rd_drp     <= rd_drp_reg;
wr_drp     <= wr_drp_reg;
not_kill   <= not(kill_reg);

process(clk)
begin
if rising_edge(clk) then     
  if(reset='1') then
    state_reg   <=resetstate;
    holds_reg   <=(others => '0');
    DI_reg      <=(others => '0');
    Address_reg <=(others => '0');
    wr_drp_reg  <='0';
    done_reg    <='0';
    kill_reg    <='0';
  elsif((lock0='1' or lock1='1' or lock2='1' or lock3='1')  and (not_kill='1')) then
    case state_reg is

      when resetstate =>
      state_reg <= load_addr_agc;
      done_reg  <= '0';
      holds_reg <= (others => '0');
      
      --AGC LOOP--/
      
      when load_addr_agc =>
      Address_reg  <= "000011101";
      state_reg    <= rd_drp_agc;
      
      when rd_drp_agc =>                    -- Start Read Sequence Wait for DRPRDY
      rd_drp_reg   <= '1';
      state_reg    <= wait_drprdy_agc;
      
      when wait_drprdy_agc =>                     --  Wait for DRPRDY
        if(ready='1') then
      store_di0   <= di0;
      state_reg       <= mod_drp_agc;
        else 
      state_reg<=wait_drprdy_agc;
        end if;
      
      when mod_drp_agc =>
      rd_drp_reg   <= '0';
      
      if ((lock0='1' and lock1='0' and lock2='0' and lock3='0'))then
      store_di0(15 downto 12) <= "0110";      --/ 64X
      state_reg                   <= load_drp_agc;
      elsif (lock1='1' and lock2='0' and lock3='0') then
      store_di0(15 downto 12) <= "0100";      --/ 16X
      state_reg                   <= load_drp_agc;
      elsif(lock2='1' and lock3='0') then
      store_di0(15 downto 12) <= "0010";     -- 4X
      state_reg                   <= load_drp_agc;
      elsif (lock3='1') then
      store_di0(15 downto 12) <= "0000";   --/ 1X
      state_reg                   <= load_drp_agc;
      end if;

      when load_drp_agc =>
      state_reg       <= pulse_wr_agc;
      DI_reg          <= store_di0;
      
      when pulse_wr_agc =>
      wr_drp_reg   <= '1';
      state_reg    <= wait_drp_dy_agc;
      
      when wait_drp_dy_agc =>
      if(ready='1') then
      wr_drp_reg      <= '0';
      DI_reg          <= store_di0;
      state_reg       <= lock_agc;
      end if;
      
      when lock_agc =>
      if(done_reg='1') then
      state_reg <= endstate;
      elsif(lock0='1' and lock1='1') then
      state_reg  <= mod_drp_agc;
      elsif(lock1='1' and lock2='0') then
      state_reg  <= mod_drp_agc;
      elsif(lock2='1' and lock3='0') then
      state_reg  <= mod_drp_agc;
      elsif(lock3='1') then
      state_reg  <= mod_drp_agc;
      done_reg   <= '1';
      else 
      state_reg  <= lock_agc;
      end if;
      
      
      when endstate =>
      holds_reg    <= "1011";
      DI_reg       <= (others => '0');
      Address_reg  <= (others => '0');
      wr_drp_reg   <= '0';
      rd_drp_reg   <= '0';
      kill_reg     <= done_reg;
                            
      when others => state_reg <= "XXXX";
    end case;

end if;
end if;
end process;
end drp_wr_fsm_beh;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity lock_detect is
generic(
  usr_clk : integer range 0 to 4095 :=150
);
port(  
  lock0,lock1,lock2,lock3,start  : out std_logic;
  count_lock_out                 : in std_logic_vector(31 downto 0);
  dclk,reset                     : in std_logic
);
end lock_detect;

architecture lock_detect_beh of lock_detect is

--signal lock0_reg,lock1_reg,lock2_reg,lock3_reg : std_logic := '0';

begin
  
process(dclk)
begin
if rising_edge(dclk) then    
  if(reset ='1') then
    lock0  <=  '0';
    lock1  <=  '0';
    lock2  <=  '0';
    lock3  <=  '0';
    start  <=  '0';  
  else
    start  <=  '1';
    if(count_lock_out=X"0000000A") then
      lock0 <= '1';
    elsif(UNSIGNED(count_lock_out)=usr_clk*40) then
      lock1 <= '1';
    elsif  (UNSIGNED(count_lock_out)=160*usr_clk) then
      lock2 <= '1'; 
    elsif  (UNSIGNED(count_lock_out)=640*usr_clk) then
      lock3 <= '1';
      start <= '0';
    end if;
  end if;
 end if;
end process;

end lock_detect_beh;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.NUMERIC_STD.ALL;

entity counter is
port (
reset,start,stop,dclk : in std_logic;
count_lock_out : out std_logic_vector(31 downto 0)
);
end counter;

architecture counter_beh of counter is

signal count_lock_out_reg : std_logic_vector(31 downto 0) := (others=>'0');

begin

count_lock_out <= count_lock_out_reg;

process(dclk)
begin 
if rising_edge(dclk) then    
  if(reset='1' or stop='1') then
    count_lock_out_reg <= (others=>'0');
  elsif (start='1') then
    count_lock_out_reg <= count_lock_out_reg + 1;
  else
    count_lock_out_reg <= (others=>'0');
  end if;
end if;
end process;

end counter_beh;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.NUMERIC_STD.ALL;

entity hola_kin7_gtx_agc_loop_fsm is
generic(
  usr_clk : integer range 0 to 4095 :=150
);
port (

DCLK,reset,DRDY     : in std_logic;
D0                  : in STD_LOGIC_VECTOR(15 downto 0);
DI                  : out STD_LOGIC_VECTOR(15 downto 0);
holds               : out STD_LOGIC_VECTOR(3 downto 0);
DWE,DEN             : out std_logic;
DADDR               : out STD_LOGIC_VECTOR(8 downto 0);
kill                : out std_logic;

-- input[7:0] usr_clk,
state               :  out STD_LOGIC_VECTOR(3 downto 0);
count_lock_out      :  out STD_LOGIC_VECTOR(31 downto 0);
lock0,lock1,lock2,lock3 : out std_logic
);
end hola_kin7_gtx_agc_loop_fsm;

architecture Behavioral of hola_kin7_gtx_agc_loop_fsm is

component drp_wr_fsm 
port (
lock0,lock1,lock2,lock3,clk,reset,ready   : in std_logic;
di0                                       : in STD_LOGIC_VECTOR(15 downto 0);
holds                                     : out STD_LOGIC_VECTOR(3 downto 0);
DI                                        : out STD_LOGIC_VECTOR(15 downto 0);
Address                                   : out STD_LOGIC_VECTOR(8 downto 0);
state                                     : out STD_LOGIC_VECTOR(3 downto 0);
done                                      : out std_logic;
kill                                      : out std_logic;
rd_drp                                    : out std_logic;
wr_drp                                    : out std_logic
);
end component;

component lock_detect
generic(
  usr_clk : integer range 0 to 4095 :=150
);
port(  
  lock0,lock1,lock2,lock3,start  : out std_logic;
  count_lock_out                 : in std_logic_vector(31 downto 0);
  dclk,reset                     : in std_logic
);
end component;

component counter
port (
reset,start,stop,dclk : in std_logic;
count_lock_out : out std_logic_vector(31 downto 0)
);
end component;

signal rd_drp : std_logic;
signal wr_drp : std_logic;
signal lock0_reg,lock1_reg,lock2_reg,lock3_reg,start_reg,done_reg : std_logic;
signal count_lock_out_reg : std_logic_vector(31 downto 0);

begin

count_lock_out <= count_lock_out_reg;
DWE   <= wr_drp;
DEN   <= rd_drp or wr_drp;
lock0 <= lock0_reg;
lock1 <= lock1_reg;
lock2 <= lock2_reg;
lock3 <= lock3_reg;

I1 : drp_wr_fsm 
port map (
lock0       =>   lock0_reg,
lock1       =>   lock1_reg,
lock2       =>   lock2_reg,
lock3       =>   lock3_reg,
clk         =>   DCLK,
reset       =>   reset,
ready       =>   DRDY,
holds       =>   holds,
done        =>   done_reg,
kill        =>   kill,
state       =>   state,
DI          =>   DI,
di0         =>   D0,
Address     =>   DADDR,
rd_drp      =>   rd_drp,
wr_drp      =>   wr_drp
);

I2 : lock_detect 
generic map (
  usr_clk => usr_clk
) 
port map ( 
start             =>  start_reg,
count_lock_out    =>  count_lock_out_reg,
dclk              =>  DCLK,
reset             =>  reset,
lock0             =>  lock0_reg,
lock1             =>  lock1_reg,
lock2             =>  lock2_reg,
lock3             =>  lock3_reg
);

I3 : counter 
port map (
dclk              =>  DCLK,
reset             =>  reset,
count_lock_out    =>  count_lock_out_reg,
start             =>  start_reg,
stop              =>  done_reg
);

end Behavioral;


