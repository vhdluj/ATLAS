`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Cz0ATyGAKzjDWjvv91NpKN/mPQyCZwjQS2DoSkZIZqEBuKINiDFaI7lAnirhiywoAHcRhiTAoHBj
3FT78bTeMQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ivOES8cu99hiNLTSHoiiiUeUQKx8vN6fgbbxtnrGa8v7e7CZ7eayAItDFvLXG6w7wbPBCOzzvjmM
tAbtGCVHcAgKULPu3afcHy0YiB5KOqCgNe6LWu6yme6eQkcc4BTJxuYAH/N+NlYHMBtBNeTmYbYC
bdF1hPQD500x/10n3jg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GmZ230kw+kh7TAqLsTElI0uFKeUHAkEXy6+VMt5CYbApdcGCeQyxl2zRHbc1I5wO0QJ88V3OHrA8
BZoSb2pp07v5kLpV2XFAcOk1BE+HML/Pzek6iUXFoj0SQjjk/eWIolmZi71ywPXBnzAp6KdOULHU
RqSE0MdIIg5rR9mG7lwXvArloTr7U4jUsQKH6+zlNJ5b1ySNF6h18nspdjzRAXBVdgd+9w/BwuMG
GTbJQt3n/Pm2XJEuheHB/ImfWJniiMHSg8jPUFzeV4z29Pa9WK06MFmO3PhrcFEhE++Tk93PxQYl
tylmhwBINxlj4qALgbkq3DeMVVqIqg5ZQTtjCA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GdrDSyVLzmUVnm/k3zQ7WbGQuaqzd0UwbocMfEtQigg/aOheHjBKRglQK+CzuOtPGhZciZgVR9S8
ORLrtPcEgDKbvM7hCDD4pczW4dmcUeMYR6QLCEVDmJUM5uPBFqrTmHUaziwSink/iGlDO/zmODEj
ViR1fYO0cP0neZeJ1CI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bIDLkqIvOvVES271QPdrP077UFYJexlS4d+ZAerBaZyCqB2UYlTvr2qpblOKwJP7wlrbzPRUAlMz
e7S4LSWq54iZn04sMS8G6Ybauu7q1iWct8nFqZFDYeQOAlEAZ3UDmcbfjA6/2FlMg78h/bUC0CHs
934K58IbtU7bHiegON1Krs85eYxlcjx2aisezOkv8yh2RaEiQ2ZEnhU3LCaIIKkR6zFitEF/bVck
nKDDiWegiglpNG6LE4zoZpEOlSYxkXWzxUzdCPDB6POib1TOcZj47qcbTcs54uzkwWmqKyaFnTlX
HYOkD6O9Dohaol7N6QxsWTEHYBZaxW4SxOs2dw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19568)
`protect data_block
twZE4hQRmTbEX3S1sEKEkvWlFoiAoMlW/VkHSDf7VkMH3lr/tVvCouYMVXkmtNkHJT+yGRuQmR5U
OjP+VMUSwYJnILW1Jt+S+Leg7Z3rf2T53jgOucbVqfyrpjQGd4w70qCwYcNc5hLCXOlArcD/GPmp
2V6NQev9iaeLq2ZILMHEGf26oe58LeeB8wzX7tJDjI5NGJj0kL4xm8Dinbs4eHScD+osh3TaRFJ4
fXGKX1i6ct761wgruVTMGMkBGz+27TEQl3dqq+jnoc6/3wWrySIVaPFZcPUDrl8DVB9Dso1PJo+B
dhdkNKsB44l2hFd2KeEEiy27Ggtc+mgZmV7Na+Na8u+mhU3GvTh7SK2lygohA7/V7jQsdWU4I0VF
UtFZYhv5NmfJlLS8NJ6XXiAjGksjanSrkLRww+gmTQNb/5JPRnH/AOzV0BfQIT3KNHlfuXm8Rxmf
jHHxlxZH+W4u0jRmXOZx1y9X2efvsqsiWv/OI6W+hHg8e8CYgVL7SzatfNUwqQQJsIaZfo3JtYGk
jhKLqDjvvZ5ZveVzREBhiZvPEX+mPFglGm2ZPzjK0cJChilcs0f1hhqaMnBXkkPKnWq/1pcWAJji
TagJskKR8lx5K54YLhqfp/TRyoxvV4oWTVA1QERG+WiuQmiNZOelsqUd2De+IaphH/iWgwwAiXcq
GVjuOf3zg6ep8pEYAL8vxy3zrX2Elfqhm7MkwEp8ZcfQQd6GpnNokYeVh12Y6THzZBHU1TFRq1/f
8QpkJFqaKxxQpnlolMKN+OeRCccYYnCLhwnMfODBzODcy9Swktr4htpjsPU1nachthpZyisuaX6G
db/6pooJ6SJCojKTKJA6n5Afl/qCAQw1uPCSjjSYuAXQiROXxxHfwzS+sz++FpIwtz+MfyXH7orn
A8VyOrrgnfklGmc+7u7rthsiYqyMCBgc82Url5ndmlx3n5m4FhAsyAXSZ1Dw52VRrNGzqYj9O8P7
uKPcZZ4xsVCUwUCd6x7jZdx0UgTrQWwHimJAVx+dj4pUXHWg6QeBoPu3poYKogGoNXuiqoPq6Lr4
R4G0CNloDplyVxhqLyXMOvOMGNDUa8RDfF4QDfxIupeXyjvnGzI4dPoSYw8rStNiuiw7ms2w5cnW
cI9g3EEhNwuQH6ofWm/oXUI72ZqMCx4xo+ARiUcJ7SeE4KEIMqhXTCgB1vD4YKI8usxFep+0w/0p
OWYPu0LS+oxxA41DGUFpR5gBL++DKSH68mY5rhIfhV/fC+Q4JzwRjNbT9+GipqtMcYcvMF971RTF
/KI0VsXsVlZwWInN4ngtAgZpu+rjDI26w5HoVQKlEnMKoGanCTcdmKTy1qfR93Xpyl4yE2+wnBgJ
wy5V1ykC2+UZZI/ExWOC/KMnYf4ztulEZKgdJXfDqaC3F0r3I/Ad7jOpiehDX/RVShg1thO6asEn
7CShSrYfaUhG7zHde+GrFdujIERt7KiIJQJoqLAild18DTUZz54yridVUFTj5LlYDUv+ikVuAuGT
iK7obg2yvPmG+SlgTcaXAou8Ag9+AavpY8OhtVDayvWOejDG9/GrBbd0h8zvQO+/9sm+p85BDC1o
H6o/dlT7JsTPJLeZY+S7fqjaWFj3B4sDcQy8zR0yHHckwX/lfVrKMJbIuGSS7HRVfph7ieqL0IdE
NSpkniAi0IAvEcupcKSwC3DnFF89xM7JCD0Dx4EA/g2IOq0sp20U95DkC1+PqVC/EUtcS3qV8/BV
zwPV/q4AAH3APWB/ibbzPYez82WnlX9YMV3ZuBRntuyD5XvdGT1FOGdZ4UvSCTO552f6/cuxnCR9
jexHqhkfCdLseOAYYfqCf6YHLwEzhSVmNuJHNdqZAxXYZshBnnCPHeF8Ndc6+Mfk2n54Vo5xamYW
saTdl2Eos/ROfYCsQFXZPAeBvccCXwEVsXKdMHX6eRuilsZgFdOXFYODFA/dvP+jCYs2lk2m3qJt
SFVWjqRPAkpv9a19ux1ZBUwmnIK31/yUEdfSd5FSXLKORSCPYdmvNU+YoJnLgmGCejJDRAkSmojD
Hk7bse4K6d6mDL7hXO3X+gPS4iBQNfa9hUiawLQ4EkScQs7eJ46LVbBHQ5WlodWbiTpQGyoAy/2Q
BZsvtXdHeg0aajDtLST/DnD8YcPVLy9fZ4awo4cHubQuoPvaf2zhH7XTpVfXaYWOUFrDmfKYnHU6
w2NifHChoiYtZmH/QD6ZBu35qyv4YSzOIXdKPEChAHQi3aPwpYTlzY4jqqq9sxc+YcqLKHcUtm00
hg60dq1ViTQKMFOeTZa/aLIfW1BQDr9IrOIdjxZjOruM00IIF8YYe012zdqhk21PLL8BGkpPBPQ/
Uqe1KGQAKYfyWXSWPDiEPpdiwGYDYbGwIchekJjgd9OIfglo8GxSM9Mf49WnyE28zHQveZHCwnRt
J1UB3l8w5QgKYUWQFgYli3rNVTCepRQCZ1d7QeR7oifTS/TbnDfWV0a/QZX+m1fL9+vEmG7e/aMs
OcwDAB+RLIKGhJBU85Ty/9FHsQtCZ9Ma3qZZVS8YdkPj8l/hw9Wj4qEQibiFfdKP5k6odE6w3O4I
KNg+6E36Q7JN+enmzCOB4FMvq3b3dcrBQ7cUAkE3aGoO0pZ07zAYIFLK2AfJcQl5HXminoiz56ha
ofWKo9VXi9AYuPqoN9xg1Qp7Njb42BOvuafTwf/Zg8GV7AOVYw+BOVGfaq1n1Bv00NwbrY59jydf
aeK3zPwPoOKIn4/NKHvfFExFE5eZWjNy/Mz00854NshopXoBceAwW8ooc3bTW7fv5Kg+jBY8s1uH
WRFbXsl1CwrjuICVUBPFaNp1M1geTfjyvgNArKx7YFcu5DLBw9xG1YU0ICa+u39H52iXArAC0s9O
7hRdZOHf4wXZNTwjukq80HLz0RR+UCCrRzHMzbcwBMpKnIzvVN5u+BsXbQXpol8fw/kEu7dQHIYk
OEKiC/lj71iojdSnQA2RZOpDNHyPIZgjNvbHgoRTp2daomLWav7e/0RhAl5qvXU+MdrjiXTt45ye
XA6InaLl7Aci2xFDR4U2/47s7Cf877kxQclnJ1kVWTjwVET1WyHaJc8MVUw+x6R2t8CAu1IEwfrU
qP1SOmiFpyeHcwUTzu9sD0TsMFitz1vr3D7oDoFMGbFOibXXYxkibWeuGoWUUgDoZvOHci5HdTAM
m6kzOGMps03Jg5Zqh0nagghnJdiGHu9qQKouzi0rME/HVLvVXYfIoz7OUIDlp8bxDPnokOBTPvPv
ukKdBzuNeMWCxkUFmH7Tf0r9SSns7t3OSjQE2p0cMX8MnnOHn6kGk6Z3jM8LOfosAUCnrc/Dzs/X
Tbc4cRLn1oRlI8QsoVNqkvLf5YyAZCSLrIwP/U6FNxFba/5F6E8Fr2y2HBpX5gO8KhUml0JTNRpX
sWeGokc6tRRYFSbDQJ8pZRBFj6ud15EUrXyrabI3gypABa/dtti9KbKlFE06judaMYujY303Qhmb
WPVBRYiZbOW6KasK2yAUmZFjcYu3TPlvaxmR1s6h1kJe44COGUD9isRkt6SKS8l5+tDSUzGS4q8D
i29InMaWMKIwosSUdKTbEzh9hdrdb516eaik6lrKVrGupbBVV3YLNSaZNGLuF2vaT73IR8J/u5yx
vQavuRsi3II9ROKicTZM2i81ROAwtjLJOo4voS322ltToUxRYPHeJ26s0913Jagp5DXyJE2bNOkl
zNEgPO78JwcFVxgnYX6zDvz3xg2OA3T9g7q9tKS1hu8Oszuin66h6N7fMQCQzATJlAZ5TcKSNHkR
kBA+NvNFyLuaD1JqnZZN1Ccswe1mSO4NDG57kzQ8tkyVGmjgwa5dJMJaoQAht3XV3gznsK4iZAwB
qMSgBW1wWUovHhVIDzeoRj8zc4Mm3EmaEQnMoOkfiSG0dLD/CeGmyzcX6Qdnat/SK0diq2LJ1rFm
0onRWHuZ8v3g+Wj54K/w5aDh/MQ9Q4q3+IFk0onk/gFaCPzp2UY2Z+ByuCc+TWBsDzha1Wbk39rD
4r3Br5IEtar693uXJ0q4DseA2bPrFRxJeklgjWvebEepiy413+jkX9VxGRmtHofHtgH0dL74LKXQ
6PiK0O9Y/A08HgrzE40wMfAEnnD6fE3GT7iPfXvEbSGWereEbAPT5Sa1jRnt9KqN95LBcmMnncHy
B5BgWIIN7vWQjTH7turS2OKJFC6pWxLC/jIntAKWUw44qCu4ZWB8EuH08h7k4zk3F1OENEfF9kbg
oQFzZS2b3vTuzPWDOiurfzAoCKOXYDpNj10NYU53L4neTIzqq5CKZKr7u8ZRHcBGxypLapFzqEh0
e45aWmEnEM7Vhpm2/+4+cpF7phExo9+8AQL4NCk8673mVyPnRRnwNc87HH7FVFt9WUIOVpUqFBcr
8MnkVkLZ4bSnawxgbdHqBoc46oqEecooUa6g7to54tt38s7GBOXjws5zt5hp81aQn+2BgKCZbYUp
K/UrU/E8GmO4WG3s7FQXJwolM56ZoKWdeibfs+yGAn3B3HfAvv5KnxSo7tULS2+FS3z9t1ZjcBWl
5uW4WTNUwjMcnAssogwGs1IFnlwRpA4g90nMOYL1VfADDDhNoCskYyzHHRTE7vQylRXPGCvYEmjV
tHF9dUSkm5ihth+aPw3ZSG/PYuVJ+jWtitJDEy3sXl407+SV4KkV0ghQzDyhctSKc/7ZZ8fd8NRM
HOLpgli4kRVbEqzSJJjCNdJUNaqUmyYThsGh5l+iGoQ3tAr5s1iHdVfMw8Jr5MzirDzG+hso3UyE
HO0H191LzmS4JXtVECmERBoyQzlMsTzJZkJR1FCuxVSV0ZoIzetcxKeaUX9SusBiZRCRk+Z9FHU4
Km/MF4wH4LINAIr4KSrLx+/ySVRhb2dHKF4fJGNGwbPb23fytnhcNy2ZDtoadjMAG07aKGkbCzuz
ZpDZqyDQ+6/4kmnHqrYQ59TXJRcPYIVEgeyiuLPH4MlDpgnuZ0GTR7QuEq+zbN2JX5m8KT8wpYag
/9T2tMCH6SwhJ5oLEUX+QP4xyGeInM6G+3kSg9z61u8iBRgeZX8OKvqN9fV6sbXk67/4S67tuEKW
LcDerKEEZBzPCNTkFFKBYRSYWQe6of02Iqks8mt4N/W9VTItUrU05JB3K/UkGP9u+Nrt/k6s4UL0
31CJc7D+kQay4P3o3vac3AJ4dlZs65hqBOU0+FwOnu95Nf4Fzxs94QUK9XqjRbwZ3fgMasHfVP5D
hJboF7D597oYeyw78tmvdeeBqN+nd9IVW4l6plaKdFkD/1gtZw5POXIlgTF8pTWscAaszSh/Y/rA
bQYaw5/2y3ZeC+gpwrGzbLR8WDW/aT6sYQNA16rq0POXDlUwkQZxC/CGQopHWITW6XNyR44HfYNn
BbxxfxS1YBhWgIwcNY/P69CLHvYSkTkeKIzwdHSCoa/LIOX0/1RepbzuH+zn8Sjb62Vxa4CMVGLx
NuEc7iQrS3Br2YQVQNOsHhkU7iQ/x7VbKkb9n1KUdcADEVw1fJzpPQd+v/hSF4bAl/DRnJKBBnEN
KV/a2pPc3BCG+IgIlcXonH9lVjpJrWlVHr3OllpwDGxlAnQN1qPbHW4V1waySYprDPQ3YIcwhkTr
5Zy19SCo2e2ieeiRIwZtl5sO83ei37ntR92uLnmMl1hdEW9W+VaYH3K8tNJC0aQkCeQxl2MmkWlA
V9RAwf2DDOSfSWd/zV/7HO6/RHSoFOvIE5WD9GG3x224vXiuAE+LXI3Koizz0FgyrrQUgPQ9BrVS
kT137gio3vcka+WDbwgTp039bIjJZIu17Oj0Tol8+W7d4mzKLaSTYvBfM1yvyoS3licqkQO0kfUl
2uErchGOmBdozTX6AEMkW8oEL1e6+oGm9zlyynilmXid7MsmrEGsppJ7aShcYsBsnHM+udP6eZRe
XpyHjaek5aFC6ufBwU2b59oqWk6XsdB3Ntuak3OT8rfoSJoFgxJ/ggYNzimj5lxizceLRAIL1x81
x6pChqRvT4ENghbf1k7cmSngDE1dUKAUDYdmEovAwFBYoepkcZJNh1LOddtNcAnhNFt4oo8JGEbL
J91lsm+Rbg52o2YUfrez+KPUNvOhBgUUncBVVnBhLB3LAL6yhyr1jvAT0HP1L9WHoy+zFyBoMNQG
yXSepR6clTcAHjiZFtMpUvt9U9+7tHIL2T3sRTHbSEveimjWzw7IiwpYgUX2gm8SA7z8dkmMGem1
KQAAmFPmyAWJFAXa787P+SAN76oVQ16Dx+KbDyjQBwAaZFjAK61U7+W5Cv3PssqvZkUKkH7XNj8w
nnQtnInRbmFxCkW8I7aanJw1gTWdw2n+U+1LiQD/dT78KT5HlGc6sowz3msdQ7QwaU2NPSRLyJNr
f99Sta8Fq/VDrMkfnlHpZRULHlafMt6nYeZGAPvssUMxGtW1RV03jLHUx7ZbD/TTf/cMNaClsV3W
AEj9fgIzDfUcf7KpriQM1PFflRvx8PzaxF1SRj4A9EoLab7qfSIECSc2SA3OAWMr8kEFSehjdOMz
Qdcpsk35BE2sKJKfkxcS7wXCrH35UbeUUMREr9+WsKhjhKG3kRT7y4mbNtstCgvgqbs/Yv7yfnI+
NRsgMvuu09o3u2CQ2JQxXc6Ib9F+pAPEWugl3GBVcjP7kDLS93oGTPChZZVno19T1Yzg78vUJpkY
g6HNIvcEPsaq3745rlbb4ir7sZiIgYM7O91lyVQ/uz9D00KWqWSEFXvqYFo+YiuhJIGC6W1mlZz0
lbcoC+JcBKc3nQViE3QynTDZ9sLPYRCqZRAUl9shJaLsjXHA00KTMvV5P6fPjV6TIP7uKIKgeSpE
6ugPqli2bqdbh4xnXIIvdXXeCwsIztDJM75qOvBrfikM3vw0gh6m+T6tueJkl/EHM3JvZsSDTPc7
K41myLDG+10vifwyOs3n2FgW0Ysawpc8J09eIQLwkBX8b2Ln7qWJxe4uWQZD2bhIx2BNqTKUrQ1B
agoer7fmRQniSkgniy9Unk60Wifua2YqPlIDBVFHIo2xeaGSBV1FF2C0uS2zw2LJZx5jWnaXh212
AxC6KrLMZ8Z8nGop69OsZGzf6CVmcfIcsFwcujgO0dJBnyKPgFu1JhrlXbIqSZKxJYGEvdpT6xze
+uTpZnwz8NrMLSOcIMQVNbYbaAFnKlVO9djVTJ6I0SmOYjM5AbRoznxMpg8kgsIL1MNJUStK1GuA
SYxDSrffEdGVdv0CDxJ0bfaQMGXS+vBIo8ZnaYlXoHfLza/2fdsMy/CRBAXvZ/kxLW5u4kr2ldWb
vErFyX58reB1852b5h1HDO6SzpdlPYK2Ff7fGGxVdyVbU09GbRWrLela+l9+ej0omDA4NdV/70T+
wal4EGW4KL3rbaNZMxAWPJQPwZLzUVWnNerkbSZy/5OsIigV4ZkGaLKskeQyPExCTm79hGUaxwjh
B0dlp5DqZ9zF+lhuYHoT6vEMBwqag+zt3HOcdwtkLX4SsovEsp2ByWZb0h7KGsxF9Hk/1pXWV4Ra
boZXB+E18IzkWjgmnz+2IrYtd+67kXCoUgk4ez9qxV45/rv9cZlPEN1GZ5jGPSUY2iEq6EtNa92L
SrHMu2mw6+PS9Yl9MdNySfLae6uPJQVL6yKonHCmhE79tdj4ihSMHmGuD9FYVHbZIegzqMesoFts
DEE4+ygeSu+yDXz4D24KTDl4AaZ8jVZxM7+tbKA6QHxuJhgDJ9b4O7RtBWhAnhGv4Va0Zv51bZFt
251WzWdIzfI6hrkIIZGbs5qOOA/ULoQXRMRO45k9HzzMQuM59Z+zF1u9AFF0C86zBe6pglVxSSHg
YG25MT0kEMuQySi/BadUNaCo1v7ix4a+F4169yrOZoriOzOgfIlaS9uG9RMBFHs/PO5e5O2whkw7
DfDsUxwHlBIs8JYDHlj3xTns+kTx4+WSVeUJzA7/fJi3xzzwLVawv19QDgi5GjNAgg9E1o+RpMCh
QAKXDvNqNgB0RNwWNYImwrIcOe2bjgKyM5PyQ6ADdesILfgPelEbDh+DqJVWygTlqQg7rsgZLtk/
I11a88U3K6QHIIcZZnL9V88CHLHuuSEhp3wD+P01rq+jDehZRyRLC4h1B4gizTHwTwDPMTvG84Kc
8zGcioWNxk1gYehL708lvoGBYcoQUsgc39hLdqYBAxw8HXwGuCL71kox4lkb0gYcT+DT7voogzD7
/7DGKIlwFff2Oo/sEfu/ND9jizFLS9aRkOCYm5F5Re1o7s1Rj4VmezSfz+E9i+gXWahce7Jm1U6i
XShywa4QXc4pTCSb3LkjscuDJGYEEA7akXee1zjc2YTnk9HZn9g1aa057msM7FOm7rAnS+cD9KF7
boI3l3wDX6xAAg3CD15QZ4SWtjy+NBtGzdlgTbqa5pegQoMgvptmksxxeaL2ERWgqTyW85NbNMzx
1/0PZSu2SxVHFYqoKLMTJ6wWO/Z4Ni/UhDChE83X41m7nAXJXP2V1J7tUlvuiROc1oNF/9X+GpwS
d3+EfcREPlJ+ef70ztyJBmHas1lqg6Bht2h9U+CLg3TLjOqeqnWmnGlRNMuDD+EaJmOQNNuWXHNw
LoF2E3G6JZs9az3tpboec1ZDTEhEE8sOwpZt/KW4tpMV4owTiiw/oDuxFtyTJRgKT7a7skxNYx1u
Uawmtvk6Cw9+z8f4ntoXUYb8tH2ssw+gYu0+LhlVuSsy7EEGeVjqvTFXiKz49HtL1pR7hi9j8IHn
Q7ptgQXSsC51SbHl/AO0wGSREq8NWVZnP8zwJAVD29uGTUcPXOKW7UU5ogSVHqSXMt96p+2afQK7
FNao9xcHoOpLfAc9CKEH/GW+FMv+PWQvnR+b4o1TxFLyPvqkiH/RxXj1sIBBV40AMowDg6teZIKQ
4LqXYL4oIqF6IGv9USPa+Zw6zs93z7Zt3gVsgjHI19YygESrh9TS7T4RIyu6Ldno/HeYM/hsRZC5
6p7uoL5Ogml2DvwVi5g8Ypsk3l515TexRGwe4qrqKRgLvOzcIFVD8wHyRuNBZsBic+aV1Uc9+CVv
kc9fCanjXkOy78RBLH7HoWUC2jbiULzcFGQQtGEsaDvcGk0wJ4VTSHb+/eB1/yCf4T07tnYgZjob
767Q6/XnS+Nh0veuu740Y+b+87QeEXY1AdggcE17C7LSL5K8ptyj9tgIr2WzKt/jnYQfKzhsahQB
QpyKToNFmyxST9jDc1umM7wq1Om+WlUdsHL8+NnJ1NuCy0oot/PUMnBCuNAPK9qO5GitgzqpO/F1
BdMX1N1IQSx8sn6wj8MS9dmrDCxrpsPj9g1i5wg0LE0PIwgV1DyDUKCR4jfC0gBR24SP1iRDRJCb
PJb71LXCyQs0WEK16U7GvSYPgQmN6ehdk+hTaS4jOlpworWfy7nQra0pVLo1VPw4RbM4cZ7LcxLV
wN/bIAQD6SijCsdNtUgZ7TETDj7yPuAMPlnWrFQC5I96Z1mJOQkdFBKBQ4sR9vSoVpQHLDfxI+tX
4GfobQ62EY8cpjkPak8P+o+hH9tlCGQ7rYv4mJ0ydbd5PHanr3lcnq7ysJe6/Q7Ut8jDNe7+phIc
FLbYjeLbnTiTEF1cwKMOQ54v429o4sSjaJnkPvraRVZ+EMIEGbdQr4Ebz/Kh4b9yLuLYx4XwX+cK
FQnZF96vK5eT018DO99jI+p7VYYK93K0RMTKVYrMONiqdCa2LsAzurC7vqoLcSpVlEVl8va4MfEH
P6i5c0diiqjFNOFqQl9yubKHX+KzGVZMWidJBxzRaCOPi2N/C9my+GYSkauENeFrMSKAci2kRPl2
rC5VIbTKZicP/HsbsgiRfbFFbhxyOgiD3mJoJ/uXWDCn/lA/4wMck9cPHxkuK8XEloGbpSkXS4Xg
th10XrYux15pcdxqy2HKEQ1AnWR3BMz8YQB8zAoDBFNILWwNGdpDBFDS2xAhj9/3zF8xZSsqONcq
gtx6P8TzQDPfPyQRyziCAktX8Cp7IQl/H5ds8tlemfDJAzXWY7SspUacTp2jZqxpTOAmKA0Lu3Id
ASqH/BdD6lMupJCeO6kNeZt8hYSSh4/HqihTeC1cnWjDUBDnua3jsSWy4x8bOSrwlgchOCuBxV7X
LidwnL+lbUkQp4stWN8ebQxB/7fgl+vfisAVrt3XPxepyjpdAJLx/fFuTZOh3nsTdWkwY1RDNgEP
DEPfREZYnUFpBO3DuEM+NbX2aXgY4go1Uvdw2M2T1VMfo3uwtKYJY1+g7bZZzCAEBtHlDi39y2Oz
sJtzgVn29K0KFrZfpE/elxOnKd+VTW0qmW8V8n4m1KBVmZRAde4bF5uvtdMM31mVGBNGNGegvkba
LuIqmUUv7MQzJiWQIgssKvYeD9WivNSGHtLg/cQP+TCw9IFpi45QKhHaVWyd/JaxRi0mffkKYemJ
I3ehXX2FlEjKg26KE4ndvooH2yPXarXTR0cfagZixR442DJTpegg748qgtMKGfVo94CHssxgTLL7
A/kX7q+7qFPs5aXecQNT5UcQv6cTiO9qXfREA5tjFv2pD13wwaeg8EIUGCFnld1kLH5xz0Xi3v3o
ZSL5LdbyZoLbmJkcUozcBBT6ip3qsw3Ly1ENfY2MfcfSuXeaL09EbD/68HNUf6l9MRi7T9raScIn
/RQ+w3eOXbzIsl8ks2rKe0RsFFQLbeM0cK/n7Jylv/Myk2HyYJYWCEevY9AComiJ0n0lWIZzDSPz
qPYQnXiAFof8+yD24vExxU2EEmV74OudkJkyczQaHpcOldmYLo6cLqqEc/A/RWAouWlPg+U7Oa7S
0z74ZDQcy6JWC3jE36TBkNr4CuzG9Vw1MyuAvoBjxT34F1ZhO5NLIrTZNPBJjMPWG14VQYwgWRsB
CZTpvxbkd4tprwPiYM0AaC7mvpj2HR0MusqhZDHwXbc3vx5su6XhRyM+SM071P2VMPHEQD11blcf
Ca/YBnM9UR8CTKduOfVlf2lJVx+kR8WHbGmMay1OrgcQLCvFRqT8WKcY2n+GK7oOea6FsmADsGEW
1w71UpMHgl2se3GLjxAhKvjDkznEJvo91wil65Db+wlueLEymN7fTynqnHbq6nyH1oN+jwRd1iwv
7CcSFWovxWQZ+GdyHqMrSa9uFDgbnjVaWGhEq510R77BJNaZYTAQ+x2H0NJ+moHOXbSZu9RKg/3B
V/2whcNqD4be9T2P1Xt6WkfEbVxAkK87FltFgn7T9nBkKjzfdhTXI/sUav5eGo9rnekgEjRd2fGM
5RVmiBvblPIHPrtg36gcRESf6893UwaLYSiKHQriUZXLxrBbABF3S8f2/UgZQZk1Y1KrOYn4vNLt
hNYlSqErQ5FLwxlaE4WzSmpcqyPl5VW2qXRvGF+oiYcteLZXfmllH7cH/RZYhnrKjmKoy7TkuWGG
LiiXpHDkdbhVBri0T6XyK/tgm3P0FKe/qb8/LVjHrvtRhOUKPfWRt29kINDNF1cEy24R45A6gOms
pVhcHn4OPDr7H8rETBYI9zhMJ75rEjsFJLFkzbJKTnTtkDtcXJXMgnbFKKYNJH3xJnA0zhQOc+U1
NI67JEJe9yfNjYe0SnfbwcbKYM6lw87r4jrykXIRepXho9lVWzlmz1UFxRX0Y7xlzCcTY/bwopSG
trA9e0DbcvhIT3r8RV2TScSskrLLw+8yltcjf5ogAIj2xvJM0f0j27Ud7JoRdr4vOuwiTMPhn6YB
77I3v4Re7pO+jlIE0/OdNlni4XT4BnKAXnYxhtjKXqN39Epa9IukSOsPRWXVmKf790jMzSMamaVz
VaOpmDl4Y7cOjpbN9fnejTJhwL5C53Yjw+Q0/yk1mGmexBqbscUyxSS2wZrW23o4mTTWBUIhcNK+
y4TIb+OmuxdyPWnGR8YtLboXNlnfet8kUvzNriEehROXmyHIxEV4tVWFeMz7umixW0aBVbBon8UF
yZacoY7wvpnnK4Ycjsa5y9GcT+k/mMfMAp4rX6+mNQvtyEDgY/4OrYCr3A7L7Y3wo7ucM30jq8Bg
Tb6vF5Ovh4jabqJmkf/qdNs9+jDORKcW2egJDxcYfE2j5jPJ09A36LQZz8pIzqq35f9A5zGGZAWg
ZUQ7txrbvqnp9VNSE94IPiEUdN2t+E7oL7ONkd4NBnfGCjth8+/6f1C86idP3VakXbElmOr9CYEC
aYXmvpnbEit3fSdYweMWcvuA+QSz6MdJxtQKq1ixg/pW+1nF/k6RnBJZr2mtZVqqzqG6750ClcIJ
xqZTXFHv2xDgKr1UD7WoLoGnMR+ur0x36Q/b40vLQGV+suqVdnP6pQlrQtfk053oc1jWv8UbHI6K
sbvqMlZ59UpgnfBY8M3w65sIC5MVTrKtfxtcXvjvLosue44JytTgwPUR0YTTWVd4HDyjumStjzcl
NSctI1GXy0WPNruaWNzoPMZHyCzMbw2IAdTwOrVT1MVs86fH/P2a6QLWyhWGFfUjAflyRglfIWQz
N70OQ+ZEs/C+K/G7QvVmWbGR+uXvcVUwetoQkcUnuX8AdM18SyWWH7r+RT+nU0oEq3e/49/BbJG4
VvbdWznvKNTdKKxhQc8cjgsHsOWu3YYj7ypL+/b38P73NVLe0e3Grvhbi0Oadj1YtaeLmeOct4pW
v/XOrP1XQLeCmRuUdtWEHSK79QFelyVxEwU2RZ0ayiKG5pkEoN2oPW7+LUy/CcF+zMgZhbtVF+Hh
N2M2PNcKiCDC2lp/EC/cRxVbNOC1Uk7+QfL/cUrkqfBKMjnwFI+0ml/jgh7JkYyQE4Lvf35HJFnU
PLOLW/YO19UomzwGm3YFczHkGiLxWxoZw6yNpKR8qvKOdBf7d0K603JDcGa2yRaSi7UOW4ysE2wl
TpSxkV+jwDsPSo5slX6vo5UomzK2sFs3sVLzl+QMdMkEgdRwGfgF9UBMDWjrsx/6z3rRGmUlvQRL
YKqN5ANWgDDxSOoxhvpKgqXLojkGB+fB09X1KmQ/YtLBQnm2YodGTz7Xu9j2GVUl9r5jlulPJdWa
geugEbJJi6CpEahYInP1VjqlqnWUY3Dp++5WXKiBPhKswz8WrvAgVEkBw8ok0XTm3G0EUx+ffUNU
S1GurP+CjAqVV98/xwffWBk7GO46e6YRvqtxawbAIJc0mgOfzoCvVEvTQFTq8s7GkwEK0A2rSmLN
VxQ/TpczdlqiC1UmGrvlRcu6Oo+JhBPrU3wVkknh3HCnuYDsjLB2aXP1ndH2C3Ky85zPYIvuTHup
nHBuE7HbJHi1HR2l+EFvfSThZYo5+dV4GdnFW19G9C2Ou9kOCH4gW5nzHD9HSQ6gewP9cOVrjNvs
ImbmjHHzxVuZWGaxvCzYxBR2ivtpyurGAF/9wqSeIiWB6nLTIa8eDCtix2WtYVZzmzJnnPHodpqb
VbV3VPuXys6ktywErPwcStyYaUSyPnzR9yVD6TpMdVkwApjt7YmbKTcPIVXeKlVJuEJK5LOlD39l
LFcxd2PxAAY2t+0aEKXThPt7cs3aeJTaX78DZ/WZgQ3DqxIv6lwlqiVa8KQQn6rY961+aSoVaRnz
+817bDHfXfOovVxc5ktXWyhfecxxKU3UlwgDCmOZx+4J0Cj8TZtGaIzuERfC3vStmas5fZ69aP6d
lt3n+qtaImxvf7TpoW5zQiDH84t+ncxySSMf+0+WlnrSCit+lArAePiJrcxu3trEw4XF4Z3owv7D
QQiKHvNAk8QpW8bOv0mvPVKOtWumTiL+HhXZtzKTeA0WU80AWQeESDnxJEkeEPr/rX1w0vtGFR9P
Xu9rx4II7gELU/VRmDpe+QCr/uz7JaOOq6ssDViauXQyy2X+MqZMi3O+uubYv/DlHQa/x3nIy41q
pf852xMXIk+Jayyfilo33K/kd6NFltaKDSE1lSzvGJK7CAzn3J522E0jyqCzhMqPpWBagtkdKEdB
eUj5bfBeJIq1QV1EkU1cOgwfqScx15QZ8bTHZkN6TEt8JehjNySCEE+9N0ZAgKQtsj3hdH/H80Zz
qgd8suDbaYXABm8o3eqe3d3oNZmg+SiCCuEMDCJ0tbdNU7qlDdCxvgHxHiZYzpDhxMuf1SiJ/5rg
RArjh24iRsiZpm8P6pIYHi8sDqyIbM/GNhncBauFS56M3dODPjsULSyFKOeWmlrRmAEFn3fKbb1M
DHEmWUr4g+x7zZi8h3WuB2LK+Afx668G4hbbgvKUuR5rEQr4OETWR6Ku2vbmJPiOUiunpAml1qLl
y/Gs/SyL5u5+RSz1SpBOIFX0z8SncYLjegDriJw0egjAtDV9tfrunXZOj7B/zbKWYDEQKB8nHu/o
jiyYCZQTHwJlds30RD2IF5Z+z+X4vfjTQlr19B7hbOZz1vSk7afRM2w2FJrhZ0XdM3VwHrgzcytG
vNGQSY/+VxNvEPJMZCHzfTdO1wKdR4Qf2WaQi15UrLG2+IiflLhwIFBwqUoXuIFI79YODWVa9wow
pv+ObQUArjDKrp76+bRTafhUExxxowTrnakdgzGfmpOtY29Mk4TVSifqAfyqoU+MUSLdLsildSGa
tvkkb0XXjJ7KE7JkcaFLq93VM/uwQk0zhExgk0TFieZvZreB9wqJtRfVNFQ6GUvvn6LIyE0OmF/E
ZmQ08X0PkUFJogZlK/5julDU9v47vpab/YSEnJ9vlErbaGmLEAmbMj4BkXe980Om0isXXH1HGSLr
dR46BXV1Y3MBfuQFZ8J5k6IBvB2GyzuYjnF2/7L70mOvagRDx6KjsJ1qIPktzTQCwp75NjOISphF
t5AFDqXfFsStlonpLtdd6BH7T9XG3d9Dn87/L1bEjJAxQue/i4uKXZf/qce98GCKsb17FxTidMkR
9wGBkNtXDvmckczc+8O7vRG8DflK9IZ9dfuOVXgGDK2iZtBS37gvysgo+zcDB9/L4XZaGNIOzUd2
b+lZ67ATOkB2XUQOwf2GOYdbwhpvq2EwzMD4uGapxVK/dVqhAwDGe3S0N3PG45+pgX/5xjoF/+vO
weuNz1PdcgJdF94hzk4Cd8rbseLUVdcYkLOFROzje0moOXzVLAYrIlLlR9mOxQ6gBJwpzGqhf9ZC
/21VPHBfgA7JwAa7ehja7rfL5OBOBFyHc+U+ioqGkqe9eip91eZXFbBFReRlfOcdyNHRPVmmpLO+
2IlqW0UCaKK789bgsUZYWWJlFmIQyN/kD9ToyHAh8PtAMMTWUGXC0+ybt8wkJGGJfRnJtyFh3ees
N2e1z+q9m44JEajjZycIaQewTmMuoG0GRBVYjsAALBPweSC+ErAT58nJ7d/fZhevpUZnGidofxeV
L8xn5pGDgtBdxnau6SJopxu2PXIZmuzb14ExG18OHhqLTUCHGcBrAFGbdlyUoqcushgbl5TC2qK5
gJ+zaME51HkehFVPa1IdbwT3otWsATQ0uabtUK9SkYMeyX7Eb5OZ7xHRFIdHuNoH1ju0qtM16khB
FhjI18NwEBmcc5nsmhscuRMM5twoc6pP3JDv9BTrxpVrMZblgGjjlk7Z6moQguPsMBvTcCVnX/K4
WJDt6+HdHAi0Xmj0XyWwxvAsuoKrG9BasDieZUsnH1fmegPAoX6oyRO4ZRxgh2GCiPZ3yhlwvm/r
HuiuSNj0TZPwJF38znXU38CafYIgeiM49yljfimk9Ixe2llWK3q5s0peWiw4kxdP8q2PkzXn5EuV
gyLWY0BMGTYnTlxfLZ17RFbD1Eby2pO5Q1+gNco9ulfICuQn+6FPaMF4rODARGjc1NupgrL9ra+s
6EPqis1NBs6eiW//ORLMu5CK1dmTVOA9T2T4d8aHo9hlqHSVg9itRm/e1fCU8zUvxxHcfZA8ReaO
JYmDQOJ2f7olTqTObIMOTHOS+IM8f7NFjWmRkbKL3epv2pdToWCB4VqAxOw1K6wmBSE8gdhU/XFD
KxLC/RQYb8Fdyv+8yNBIEl6t+2u7Obxku/jowkkffJWhbdtfv2t7UpeWhBe/5eQtOROKI+gxvnaG
FbpcViM0ZixLO8uKW9XH0+tc0TdyxcexndZz9OVqjZKFVI3sN5QUa+ZEtM6sEp4SJYxOpUDWWbx9
hzP7uZfk1POILwp3ZLCXxb2WVEvVVEgypHfxX5YIRHyB6gGEjxgSyqkblce337NlUi4AxrVH1FCA
YJLUPrxBtJijCl85fOrTwq6Y6KqsD1N563LCQDWg8QFjYfvl2tYsYBtdWrtlAO0zv7iHUSP4eddQ
Tz/PY17IgsuO59UpdUppflzRSmn1u8ddSLRd+QXG47NaHJZclpJX60Rur5aeD/xRpcCM/xjJWUYp
f0baGvdXMW/a8LTX7w8Y3uSYG9VtawUvUU55xYt6fxsaKxhEiCrSbWq/t/JRbpo7g/6yxWYUHxkO
zIlhqKDuyfGZOPkx7eqfd2ODgWgwaW0wgejkRZQjMJANoq4/j9g8T6u4hoBiZ3GYdUjd7Pkb94A3
Q3+j/8DFnlAOhEX8LwMJSKIm4/kfcZ3tYpqBU6R9R1+yeu56r3bIzjjwQQXDk6KOYm9sH6eJUR/j
D/nrqbc39N42bnumOL5ky/lqsxBXMRrBi+tJZUqrHtCu0A8ZeIUygpYlvoIAK2n8OiQk3HAd+0AJ
tTvP77Y90J/Aty9ZkkTCfpwDE4vXJvcltlqQ6oLHFs77YgrVpwr2yQJi4x6Er6y1ULhvUrIL98vh
PdHxTwr5/oyKRS/SK+ZdfPBHge2tnn1l1HyMoDWtuuurwqYMLGFjkXwTxFTJ/g1eCX1WGJC4w84T
fKIgXQ1bvUjddfPgbvJiKufw9wZdCLaXwpPAN4FHDK5uuIEj3YBHSTjH2hraxQam/s8Z7a9sRUk/
4fZPZ4wnkOBfHOXORo64oTvUBZ6QQJHOjed5869lKD056t+l8TOzWBZhxdNOwaHv0Iu0qTeiRUhC
JT5J/OyWH+BquFeqFG7xtgiZcyRjhGKhB8eBee2PTt9ZpIiIXsRsEmF9+Qs5CgSlCf0Y9mlUFR8p
2CeBi2TI9/GeXKTT7dzcTRSt3imRhVd/APyzai2JArzXiU/SxnMTqfWrzUQTBU6rde1YYItC/9e5
wc/51Pmq4OzKDfjRg9hbXnTy2hu6k91Q8PvJoGOlpnlcPIqPdj8sjCDa+T1ZtxPCBR0jm3uBMRhb
0O5lCK/2WNL4tBJ+jSArZvEx51me4NrQ++XOkVyt7QOkdEhtqMxN4XZ6CvMTzdrXBEPHe1UFEwWV
RV+CO8Xxujow1QU1Br3sfTFItKaEuDL4HeJNYCUg0pnMPq+g+cKDqE993xG5CkQe/pfUVTLACXWf
BCQ4GwJet0HScGTDDrF7SF7MNWxZQWlxSEHQhNs3Pul9JVbytXyEixjY/ooSBW5ZbnLgKncUS6td
4imCoXaYmhDeS2TKKS1Ft15WgjICGDq79h2VtJBzgm/0V6HE5HLEJwRwKQSJDS1AZ6AISPEClsTp
t4jTMJHrf5eQZIGJ2IaLC/dyIN3EMuXeWTKL+FBAsl4VOy8ZU8PkldIQqJVuOJlR2aJjdIChBxDJ
iectz0pZSQzO1Sq13bqcjr8ahcqFi7tg5+SjNrT6rjVYOg43CrMH8SnQ9lT9OypYheazrzGiQUi8
rZvKlzMXrn61CeClcxzmRFY5NlxCvmxywEJtxrLA9DaaCqf8ZWP/S7fhd4lBDG9j75Q+0EmWF9Ph
idMhRdduu1roaBAlDbpu6N9zvw+7z5SIJe4tqAPUpBxYtdBcSbBH7fOBvlOIV067PVzhSgAUiTbp
yq/W1Tc0bIHj1eTqf5iEZ8tL05q75QH5r6iqSosGeS8ggxo8CXaotN0hRJqt2IMlw8h8QErl9VsA
5XGUqhDBIm1/+IOoe5EwvwPN4w/9ZhzBKWrVPMu2Yk68+1mZeoUoF7yastEEwE006Fc5lAED1e2T
8nAD7iqgILMRq0G77ilpEy5GUj0uh8yPeosXUxHcPhXG5rBMgWiw3IeSAsZu1HV+gsa9T08BsII0
G3g5DXP3UUhHIXeRtPoaIKkz7X7IbsCoyw42xdICCzS8uIlJXWXkh9jAAEa+2Miar2b81YUoq21n
zwtiXu6fA9g7pHd/XVOiwDmo+v/0qODTu9pni1Ea1ZiL1RIP06UFpFXlaf5TPbmV+fOq/4I229kH
p6gRkn/v44Oa8dyuHTLZ1DQz9v1tiycyGZMj7mGhqJTd8QrpHHAmAYrAU0JQNYOewQQRO/O957y0
+DrFUmscScwqZRNhmUU74Cf5NWX+bQLuvnIJIfwSAzISAWBLawUirPTS7V848Icnuel9fUYc+eO1
LIRo0DW3H/2YMSfl22Og9zvyAvTdAmGN7/VIik7+P7VmX31fwxIcOJJvgo3+478ptpJ6it0x6iot
f8EykkXkzfJIXgCNJaXpMTYJx2fApfXw25haFS5bIAtKtnuwhWQ6OPH3oBLCgatorIdShBk+9SfE
dIdQwxMNsQqfodeBd1rJ0qal6MlCRfso6Byb4+7URz6bbMc92fpAjhkipZojpg4Q+6XCaTWkXh0d
gORQpAhu77A6aFzek6c5ydpILb3yFr+Ay2DX9brWX+D5VTJ5lyuBLu+V3XozBI3/tzDC5q1um+yW
yqZmoJekA3N1sDDdBvGI1QHtNfm3XHdntPPNJfD/JwB+OjIFC7IAUjSOuJc+UIMxXUdGeYbvBbN7
Tee8Ji3c4A0mZu+3Ku/HZnlVBcclakJiVHOUYgwEn//Grnbs4oMT+KxntPrDF57rmYaqRJXrm0tm
KN/qN+dp9aHrKRHkR7glPv51iF5NaeT8zXfiIAX2MJHzQ2I1UTc2vUJMV71XuMni7fv3B+m8o8DV
ZQ1zkKTBkwyu9ZJOPwlNchEC8Yw6g0UdMDKGn9RKAU/o98e5cY/XimmTdjd4DpH4ywKqCUAVJhxV
2PKyBeznsgMQI0wQYtxAhyhm65yUKoFTjdhCgViYGf+ZESpokE/NiWdB215+ADLM7mPf8z5+OGEi
R0VXvX1Pk4tPMYcXEWtB9La9Y7KFkD5Bb3+euqk1k2t6zUjTciQLU7lB9uLCe12kwkFxYjyGOQCz
1UNgj19jrE/ihXqClYzDeSvvYg6cGn493O1yj/8+FN+pLgnhfFcBw6D4TjclncdiOVuVQS8YRTRI
x0kt9MzeXVD9eCes0COBMpQFc/EnYXiFLTn0n2rYcaKXN3aVOLcJoJG58Jd5ogCyQF0cdk2FuuTv
4YXdH6HrCL2R0hRg1D0g1oQMkW2WwBz+W/cgSLPezuwF777jO1eM6uSGimFWumJu2kq8tReUkOf/
rRJwlxYWWvh6i5V17LofWdoMRdy9/KqcpYjre8EUYLCwX2nq8ZQkJ+77fTVDGU8/DMsjX1gvULaU
jL041emEOqLYlgksvSYWtDwpD5U23ABuOAyBYNMw5ajM1dr5v0G01vgLYxOa2PJxbu6dG8Ee380b
yjGq6RWH7wLyiwv6HorcSsxXTAtQ+UiD+Ehho5qfFFNUxFE1HFR4HyLnl60FUe120wt+NAAfc7KZ
SHqZNyryfGCeX9eP4eROF5Bu95/kwOz8Yx7gH4L4NvFdCUIvBPxhSWOO7drGzMsFdwjAqCNq/0ma
khc9eO0Ubhxcs6voSCyE35xx20fRpuFcyGmYnKyQl/7cv51FJ+xuZ2QCEVQDIrT1VlolK64aYGRt
/7ilsYhPZASUvOmitXMpOoPIDZxDhujCmFOz7eBQaKsK+A9T+mjlVi1ya/k6+ShIKVuFFMQPi0hs
CIoAg0OhrpeYGWt8Cwid4tdd5e10JfyedueNZo4joiSBgCiO9J3bCMgAzwCOowZFwPCl5jgDNq3U
6bG5sQ7JzwLjCwSdzolzUYHf7GRg0edVcxrtaoRjZYbVRFF6uNHDDtkHruylk4xkBJKcqm3Zkter
ohUQ9hi1qYCwdhxZ6akV4anjmeJ47zQZiROzmJ/JUTkcOqv2lO2nk6YecZ157UBmkHZA1PR7JDV3
rhw3CcgOGkTe4PIkHtUSruGs7tgIqgHc4PYpY+9sEBB5x7wmMejiksjhBoEMcSY5HDxskVKPfP0I
4UHQ80PHEKkVk4wvMC7xbxqU22jLcdx0HJUs2cELmFmsXMqq0HLkWnZ0a0RVIPSf7b97EkporofH
0kXUtmGSeZlZ48HQK7S5GG6gS9YuFFy9tAZASNtIj6ueDu7KlGiyE9/tcUfcsEZXhz5NvpjuZ8+w
hFPvF2BUOmUN2c91FBpK10IoCbTVE4EwifDldKUHflxXdNWzk49705cZSfs4fMnRbwMfI84R6na4
EFN+kXSCGMiAj/1lPocb63IAktVboj6VK9M5elkcJjJlqXDfkjC9gKP0go/JGiaki8VlMHhj7JJk
4ypitJi55W7Rfs68z6p+c6gtWDLZSy/hPUphDfA7iGvcuQ2vmapRKzE2E4MNHGniqjs38UdP1y2e
YHlyWfAjYf9RdO9EF5houRVE1w7UUxsEpTc6bRMZM/44qTJ9NSebzDA+jIDXZJMosO0SzIRbVD8c
C2lw7naUZ07ttk9pPgcUvOXT0nLnfFP2gjnAv0GjlQdd7cDgR6fCjZ2LK2a+gaNPNEujq/gZdfo2
k0XCA5TzJ+ZxPFSbHGIYlQnMPYX1HDzhdbtaReYr2G3nRedYCjV2NgXmtEp5zyaQMoMwEFR9zCtY
lSfF/NDYyqv8bq/w71tBl2Pw3ohctOUwsse5+IzdBuLZY2SCTOnCSQBIJ8U2HASkdZhMsslFkCQj
qSXXtyRaecMDPHIzVsh+NqpWUfGwRfWsmssjmnYWL9gP9DCMqmDniGAAsPOymXNKPTLy5zrN/etf
0Da/e3jm0Xd+cMcUfIbo3dYxKCHgZVAYrUWbztv9uNuFU0Avu6aZSAZTAiKequ+tDeeEfMuEmqyJ
vRNv2+jYh2+qihSryfYQQ+DzwB0V9f4cgLtZkMQyu5rZoCYwW3G9TQR6wXZXWvZndhsJmzGX74y+
79frCOCI7RA6yLnwy9DwZOnpPEH3skxWtcQjBkXaNYxUihMidLXy1V8kqkG5o2LjEKaFHZl6Bt5v
o4Lb2EveXJauD+afNlKRZfsx4lMflnYDYnUza8BmWuZddZZTBahPWpm8brvrU07rhito0/SFHjwS
F9S2/T21ASXGcIv6a58zel3Io7McpOXFcFAgcjnXAC2T2+GfjukycXjIwcTiEk+QUPEMoLm3fxre
oS1eFiCnkwSd5YraHS845ucFxdTdc5FMj/rxTYav4Yv8C4SJNwUgYVQ8OKaMVOr71dPEyojHYZgj
ifAqZkxtxCJN8XXkei1Jds8VVhxUCvoTFeWm4z7Qc6nxVc7Urm+UM/cD/qb0C5UxRHBSMIgVxULu
Htw9BceTVdhXe5eINBXpsF/atFZVk9LU4qwIxpxvriz5ePg4IJug4AjhBkkkj/nF+JqM4fpZSJcj
sejMlz6Qg/HY+5VjywI0k5IEC049y/8gLL42lpSztMLwOqgzG5+lm2CmVLQHFLp9Yk6a+Hm0fMie
E8cYF97QT8FTsF/0CZqVS8j3R/le6aWL1i7qOJ5TfEpKrbXJz5NRy2qe37Q5XRzaIKmERkV3w3vc
/61cRTylRLIEehUCvjsRg6bsVhG7Zj++JtTo549znZ+LjmMu1l3KGQuDuneYupzsDQvMWVIPhPu6
hQf6js+qLGDUFjvyWyxos8CIj7LUM/rD1iQLFNrjvfHMV99mpFB7EiWR6ZPMaYUMSg72xmr+oji1
P+MApPJskLp4cW1ZJZBiCTuDvc7IKQUZGQSO2KwOo3xHOlEm9zok++3gsYQfI9ncCMdgPK8uPOb+
76Pe765/qemehFT56YB5eLD9QeRDqFmIp3xbtc+bUIzBJ3CjXc2hTBW5SBPntjZRExhjevUAOiQ1
pDp+Aom78HSg1qH0MTNWaCtlTv9Nn70N+EBZ7T1/0IKJWNl3W7Bh3xq7nLWrYcAQxeQSSEOCSnJh
7/PB6FBnA/HWQBN70ZMwBF7S0AH/j6gQAgX49duoSAi65EtL3VpRF4h9G5cGHLW8QgCU3oj0Sfbx
zv9XbUPUoZ58iEHScpG5G9ba0WM4x0+6MgDe6w5dOCwq8W5IZqwWXKDTTEZGO1UxNwwf5+wfw5pO
k+Ns2Y9O6cTl7yPvHY9usaIeFFFY3yklE05Dpz6Tk+zv/x5ZWueCcLiEdmzQF9th2PArDiFQia00
y/P9MknKq3387Ak5k9ai/vxnArKiLR8sO2BYyddeZS7s/Wi7ejSfpdPr0uJ3QrAeMfmKbbtD7tZf
dgxcJszd0Y/d9qc9PuwY5tZJbkhD1g9OTGGZK+KyxBxrsgLgLp1bN+sDuAOFxLlcqe0bBdJjn0id
dr7MSA6clPhtjnABbUsE/A3ErXb1757vzsA35FIlOQnE5I/NknguSBEBuDB0BSMBBkkavWL0Z4lo
oaSEky92bgQGpqNbHDXUSpJsCyv2UlYE1iubDPSMzGumyP0n+tikHxOonXPnax6b2zX5tknlKBHq
rEaYoL/Dy9SQ0/zuAEfC44jnMncj0iHAdtziQo2cOl1NlpsisWBF98ofOYvO9+vRXAibAh739FhT
L2j6U36OWebPhFpDPOCcAVfm4vbHM9VzzaTdqugjdBXv6EAbi7AvBLXiPA3iSBp0e1MWbPpJfukX
9oyearn/uk7hU/V/q3KaIuodFw9RKFX3CStaqg1imocemI2hU43XnON2MFwzTMBlhhUs/aMiPKtz
fNA+cWHLmAvNf4dHWsUx4e7LqOCFkMpq/YllRObR2Y9WGTJuRI7d6r4sKWsEH56FRJ9+yl0l91Gv
8rcTCw+8rHoo5i8Bjisw8J1HXuzwL/m6kA+C89wZl1RVvzq9ZkI06LkPe2aFPNp4cTfSyijVj+Te
kZ6dXlChRpNrkxlMBxwyrF8Q23J/2Xgi5qAdq8e7FTNrde5C42+Mm1iG8zMdhxaaAgKVYDzec9/o
NfPCc6JOtdCH3rmMY0FgvV1HxM9qcECacb57GtGH23XNTLG8owBzncYvGDqCS4DlhsT5pU3d9DvU
3mg6lvrrS1KwOvpIhB3MaV4a1LqpyBhA6/dp0hMfci36HLbP3Qb6bsXEwVQsuPZ8O+OaUsmzO0wS
AjQVOUChbdiCZ8mdeBhoPbonUzcZHX8ODbcZDhbavEsaK2yI+JkBphHSuhhfLo+L038CaVkOugzH
NanTpyKGLS6DG4Z1FOvliTP+DlJmv6UsYxkmtDdfpNDfDNHkGs8oviu0FmWGwSpht8/eqxopXkJv
XKgoKTChZY0k3yzbyvHjGs9PQNiMxHf6+j83HaUyvvNs71EDrFmXTNwUY1QDR9ebi6xs78nVgunm
S5siqp8g1ut/8yC66SyX9g/z/UQv6XlaDrsQMBiKbmjd4u7+RfsInZR7oR05PRimMuBk5IT2w1ez
38JfQ0cPV8jzzbp8TtAzU9zBAkOQtfFz5L0MY9MNw+1/Xi4tQ4NdlYKli+i8DHSVaGJghu9BlG2p
MCefBXkvdd/OxecK0P6fMd06ms1fHteb6VZN90uiiOPCVr2RbGEA5nlHE758doGkf0Yl6PWuX7Xc
xqR5weCqdZtGnOvX9SMO9EofzN3fmWKodp/OPnuFRJcZ0iVSWQBMtp3JSpb4Hb6kCVuVc1WCanhF
5jFqSajW4BGaWlRZ+37jhTlJqKjD/tOfZFPq32wr6ZkscM+bJ8Gb/tTLp8L8uEKO8/MpGuXY0MRi
/kkFlX2VLCOz8h2wOFCkZqFSWcEs/ZA9WPKW8VraUR9PpI3YttIOVqxu6V3peBB0PAm4ylURBmRo
gC6zhojc92mlz6h/ZafGl0wjp+BP3rCHBzzfBKSC20PdBjLWr7M/uptp5RonHXaM1sSLyZVyMst2
lb1iG38TMQylxmo2iLXp2fon+Dx1ZzUoOHe7YxAsLL6/ySWFAWoD91Ys22VcqMbBaHVEZh2T/QWY
QhcH9Rd+zFxW3eRrhOMimYBBHj9BC+F7A69IlQMxRRQvNCyLjRlsNFGy6gYesjmQ1MTn+x0YvVDo
w2UCSDAJcEfic4radbnr6KZtKFrjAOgDRvzWMLt4C4nxzbsYp0Q6mhj473D+f9no36JL/z1V/cdf
R7Hnj1X4+Jde7iFewzULvFVgpeDtFf66CJAfQApnJeWcsd7wE59Qbg6WWtkXkblMELzWB3aXOKDG
aX0lsVm7CUHV41f8VR/xmWv69ifrZZtUBp1xxNOtO2BwTY/ZBrseJbGPwMDC6Qrg3TomixHvQTTi
8pc6wWHJq2pnq+dXx5CafXjq7RTk9ACQXRou/69PaynnrJfXagLsi0+8BYSQ+gtDkbPQyY7a+1lu
EzvHJC5MorbtmZczxJAfHmW4FWFv+Izqn/oftmonQyp8+pTF2/SbZzYhh70LEa3RYPGbYa38wNNZ
YrnRwhyVN3R4cQ+HGicTssD94hlqn/DNkU5C8FbgbD+iWF2tcJaFcGlUwR0jNTPP2LijXSZ0g8L/
HXPJw7YHqNTKdaYpKmy5a18uL2AJnkLlV2s9Q8gz7zQBBUzcLATUv2U9a+2ZMs0/mQEgATE6+/Ft
8RqnqXNv2fCDb5NLGdyZWluen1En4Ex7U6dMolz+ptkWTmSuCSEq8ffk5eBtq3erR7SzNyeypCEd
DqguPdNNKs4E12sNVUr5U3fR9PRShsTYH3up+9dYXeB1smqJdxSfv5pgZ370J0nuwYBSL6BllnLq
NQuhGlCNSpQQzuQN6DykcJOae6ZShGJ/0zgqh0vVED7+FEHVNJvObSmbMDfagxSjXZp2sfqvMsYf
MtVm8Uc0P1pC+asLWsoxYeHHNjXWPQ69V22ttD/4Ixqt0B16u+MQdlQD944ABrXp1E2qwdhBEqPJ
S8/NnV02RhWRlS2CRxf7v9WTDWsasrPsvaYsWDAyv9UgRGX+h/KCWJS0VpKL+2m7Y2iAFyTrPRGJ
39Zk00ivk1K4xWrkKKeztd8Ba0entgN1j8JG+w+uRw+4XEqQuiqy+72wYNK7PbQMNKgOXPzP220/
NbwhO2VQEf/cX7Lhs2GBU+gw74MkkL3I+cjLCjp5v1dSoK0/HxqkkwxGnlgBlfp2AEX9ugYE5Q2+
Kku+wGlI4Fp+RZR2r7h13aZIdzBKax4BEQGt6fZmJXuHWWTPnjcHxisFBuPXPaBU15KwIJcxwjy4
VZfS/VDEKdEC0HNWWQkT78v5Y9gAJuFrnY/gP4BIHKk6GWHb31XyDzMlLzwtG0R4Ps0ep5qfn5xQ
W6ELSLVVAgG4m2iFC+c+Kl4XPT1yEzMPLltOIxJ2ALNtDWUS4uvIox3Fs0d++FeusuIzfeVLrxe+
a63aI6KHx2SO6wXhrJzzt/86g4SWszur/m89Gs4+rkVmoy/4r0CsZCQTSD7OOvflinqzYJReDAfC
sTsXA6yjnIARaUTRrYD4waTerhpjNq4/SILHSOFX3fsHx6hvPd19ueJDVRw55n2Lz4IpCHFcxQUc
1UHx2RJaOcTKma0/jOnjHde5mqn7PJm/hGfJBemXK+1aExMUDhtjzOzdudoyQqckNgyoUkmuS00o
MCfoZdyylKcYkAI6XBTn8h3zUo/DmJvQ47+00Ozolgnygfr16NIAVoi8lTX6xloaF+ysARiMT5aZ
qziLZ9T6sqzQwUl+fJGMG9n7yZ4Wlu5mnAgjt4ximYNJx9y7hRKzO2U8mcAmybqx+eJg7HKnnV6L
DC5vNdoxSIgMZPmL815KmJ8uSxrhr0z+q9ws0fL70+8O0oSkDmsYs0gGwi/yA2EbtpKZjBDJ0vT/
Rpbbxm9k5sMdY+RyW8OEMpQS/1jkEPSTKv65QsLsRscxwxEYaNcdBM8YkqWrYaeYLg0NEjliUsqP
VtyNEb1TxuSCZ9QGUwXlF19x/GB+hOa6t57CafF3D3e0QlmxuhCJ7mMwp3bfzzClUtEj3ebmmdOz
rkN+iw3TFxC57ZHzvXFFONaGlvH0J+rUVKD6njxYhvThyXm7SvtHwejKXPi9/iTY5ARSv9CHQrxI
ZWXhnjzkGEpixuUsqYlOF1tBIjqtJHHt3KNjSn03LVHrGX9JgE4TiVL8IF1aroH32U4ub0wZMJSK
dGI035FxvRKUqu2Cu0JvBySfRmazzIMcjH91mzssfjidpawaEMWrzwqBYU85aX3ZavgQwA65w6y1
TbiF3km6hmNCzInBFgi3gNo=
`protect end_protected
