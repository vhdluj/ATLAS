`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mSstZUXDa+xY3HqOgYFW0NX1G/O0v32WVvHeNwhH70yIj1VMeiz4urN67i6Dg0yFJBt7pPQhh/UP
xCNOimTRbg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mub3t61i84HGczBtMEWGGCYadreKOBqGj9kPUWwJUSRDfucm9oA7811GiUaa0tZgE4xJOzST3sbf
Pz+CcARN1q5N8nwBtac0pKtvs5CNiPXFsauAET4mHlNGrWVziwWm/iq7h1nIibZ2GPDcVyIxvW8E
XhpUK3Twj+ktCvcmCwI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oMCd0ttJO9NW3LLgOqJhO85ywcE9mRVxJAdqZ3CBDSUHKN2xI0Se5NJS975HTF4BIlqmqYdOC4Af
niSRn4pe2oL4Z625Wf733WSJfOOmOpYBs6Wt5LLbxajICMd3on/Z3Owcva8/DWjdd2ZF1XmJMazt
ygDgpAOJl8XrslKXAOlJHV5AHPGzpKBF0Bbak3miEn3vnzzZqHMWkRU4ZJXjmWKEzpggr4fTSLBj
VSBJbqvgNH4+vnieJsYnuW/Tbl1UsjRAxOr1086BETjN9LXFYIlytpwEyGx0iPB+5QXy6pDmqNgh
/njiyAZ1dmVUGt8fD8JJPeMG7efeKxiXtvMrIQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KGkpRkYYBC6CrqrQloFElPjv+FLasrrXHMdCaBdSYKg9a3ZUa67xOout3scZOYj7EDbM2e1g+z3d
VQCy0XHE1doHsV1FISm1WW2q0clPj/gnQZ0e8dGcqmwDQvGwnoCeHLfLF/X2n37Wx+J91F0HrxIP
rUtr8TyhZy/KtrH0Szw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A8J8O32OKfl1OLVULU1VxYuqW1+Chui3og8MVBG4ejhZqKb4RBlBN1Vf6XykJjvsOeblOEJnbP8o
mTHeY739yNUfB7cxiunuNSNMSpHeV+Jrk+0FiZosdJiFNtfFLBCdeK24low/Um5E/7r2sh0xCW/y
OZp0vFuc6F9Oqf+OBBSat2sDs1ipjWwyWVwUw9KT09LPZMM45hm4W5bGP4Ff9mYfMCvXOyoLZpQq
3Do0ZE3itmR4Y4AuRBAuxobSCq+VsL6kss9UvevvovcXH8QQ8wNk98GE6sr477dy+8y6URgWsCB+
LevrH48B6eP1jxyxpKZzpz3uo3fNoc8efFB/DA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10784)
`protect data_block
pTHtj7TIsnFHUzE+Yu8hgTkEpKf3rsekBzcjKMz1lXq3vfC7rfu9m8ODlQcm3T2Xah+Kjj6I+zX1
O1hQEAk5Uj/q8j5sGCFXyjgQqx2eNN3HQqFHdsfQOxLm2pFgM+ZXKs1zmTuuNoDQGWnZWBEne0S1
tOukzCDk1ubZokAWOoWWm/y5/Cy/FAqENuMCdaEIJ46AHjR/eS6ia9hc7tVv38251wgxfsnDj7AI
vIdMS4yQBN9hsqAv97Rak3o08xaXZX/+fkFT53D0w+pZvuboSPhMXVB1nVl9Z02/WTNEF2uaRXck
OLwCyMCLJHUknB6fniSHd0Uj+oZRez6iqINxp6n7plSIOqoiJNImheDVkHRnAZ8/6PjN63l9T2ac
CzQTa0fjdmj8aBH0QsByI1Uvzo7VygVx0DVCYfXzuCd6bqZsJg7Sh+B9+SmTyUKWyh++jQajdf3R
EzqmKVw8xXfIclRUiuQN1ATyovSiY2W0A39szF15IwcLj44pPxLv1bX3xRcaDQHdfDcql8LEi6F+
n9XMQrlkUt9dCb7bscPdaMUnhLXwkzKIsWR3X7bCfKQfLXBPQ9+6WqZabu8x9Wnv3n0u2jPZho5q
B1SAx8TXi4p3utiwLyChYRylvaLl00Qjnv1WGJrQbETrtLHUV2gvqDFLm+p9y9y0067cCkSKrL2W
I6n5QX8SiTfrQ/6fi6oFsELNRXyJJMMGe+HEtx6CJoa6Exg1cJUNRpbul1oVA99JwTCnKBAU7XA6
cn0dbO4dOIUPpCH3PtpXLAMqQbwJxF9ay/i00nZ2Yn9R2evfusGWsQR1irqgknQ/v5EHIebOQ3ak
8VyGt5nn60FbiPUnMe2cX47dw+Zq4dxWe2itBNJpXwat2eZ2OAZ5FN813qFDeogfwgjVMgj1Jilb
BHsGzfshLADRxt1X/j4BQHmiJkv+r0sfGmf7cJBhsDeLHD5faH7YMiMkU2OIgS+UGKA8BLKb3R75
VW/wmApi0LTz7xFkv05BseP+idpwB7+nk1nY2Fu6/RRG7ycrvJuzDqqjKJOSxshjp+dJH+YW1Ezq
Bp2BkpDA3O/0fwCUQzXIaRJOKXECgvq5n9bMtYASuOwKgm9D3FxdPp8HPhb6seVWixFil5tN5Fj4
y2aVC3LxJkP1wiviAY0PrupPIlB4yS9swDkUHODC4cLfcOLveTWGul9936XEwT4vOg/KY8SKz7w6
XWHu22wymc35FAyVeDwNxnNSIRYxJoEC69XIHzIOSeLOPY1i0v/m/YZhEb7knuSV7h6uz6pW1knX
0vSzqryRCzq3ecCtjFilvTzAWf/eZ/eplMWdtCbJ/hfB00LdGuGr03+gnwi+YJmmaJ3jxdbMsk3X
QL4sqODB3RPOasmFuh94/P9xjyYUrwZ/a09FRrmiGhRU5GsjKRliLGjFF1DfLvYjxyMD9FBta57I
hRI9abcoG0G3silbWDbwwdDOlDtLwi7q5cDZGqIdNBXRQmNy4Na5kqBM+Us5VKBHZn7VZemAnTZr
jzr6k3cIxDEr8rf5cphDOsHDIIX9fc/osOR7pGw7tmc/jbTZMoVR9Snw6lSeW23iBjUm91CoAG4e
IcIAKXhOddRZDKsMMm8YHHIWIJfvTpBrjS9ynB3P1IAnlw8zRNa3SDqmJX9FReY2KOEXkQy0CjT2
HqSRyubkFAtUbDt5Ub+viZl85N8DsWwdItft6bv7ODTEVIzbO+JONhT4AeskldczrNnzrvIIMWIi
7VGrUndCfnRVmxMtWiaCMOJrErWb6PCg4O0FrnWcedEdMI3LU0zg1584eTaV7ncDbYyZSxWGuPZb
r0xaIX0qaxNeq/VPfBuGLEO/61889fw4Idt8GCPiFETzEOct9ZUhjN0VmTkhwkB++Mlgt7c1b+hQ
V/e0QcDFA6BdzMWTLTN2KT1+JDuLt/nlXdwDB6Z/sGtkHeoGda3yj0bnA1EJAkzHZ+FlW1sH2VTv
W0pMNc2GQH7Fhv8xz2RlrYAncz8RZ35+VRwIu1WyYdsDvO+R/acVVWjQfSOHf8s5osEtk6uodFiY
9Du+XYS/N2CzH/NVJIOeQTzNvTuMsr0RDOmBwltJcz1HZEhQCRlzRonFVPwzvD5wo7fakyqJ53hP
JSdKF8lb43AWNUIhRtOFRTwEKXSY8Klro3gmwbM5481/Vx6iOG+19iW5sz/0xc773ghJ3nkbSWnD
uTq2ApeD5Ih+QtoV7MLaFLeTKCePg0XIlW9X0sqZmfrBMPMIfQQl6e7yPHmNTW8fT6yqflW6yV6P
UH2dtg5tUtk8cmKGHaDkmfELgyrjntEh+pH8QG4DnE0UeMLpjBCdQpV7ezjKJj83r5ppF5Je3+DH
bbuB96DhdfJ/uWo9sZ70UWAxEIpga/2Q5E4Yb2D9LfA0tMcHtHyKt4EGJ1hUKoxfOIY4q8jUWnzv
vbd81o4DfzlFPYi3gK+3FlCUP6wXmS6YgCKlO5/eRCiI6GopM7YAaapt6LbPqCbr+TKeyIFm45aG
0+9M8aUBxYPgJDVwL6lwrScB7I9bkdmsI5b4gkM3viOVe0CWMopoLo7vWFpeDSrH4T8jPWXeP1aK
GDgADIFjUm7QvKOcWgeSXC52XKHFUXP0Be6upzDW3O9zcvTgjg9mDumUa6h7Fb7XHrATQ7pii3wT
g9rh4snJzAp5pvwON1bLIx51p88c8GBOewtWzBheBqUeWlVJnlQ4KbyEdaPfjcSEodiGT/J0yXSO
YQU2vVDbx/6pn6MSA/cnnNMBRHBZouZ4/Pi/bms0ijmXt0xCFlbBi58VUAXYvI7syBJNxCoHSBox
j48rOW4K2xhafpXtBhU+Vbw4vkjpNwAkwe/Jx0LVHzEzeskRwS/jovVbd3iqlwRc/pHe8sPHe8NU
jljS15v/Glnnsdj2NEVaGRvRR7ywuS6DoubiPxBC/ckFIMTJsVUnK8UdLGB8Y0Tq+QPIX/EUeF9e
sjgylSmzaxHQKsUpbIM4EY9jYu5uVCVsUFv+FRxdkyLd5WNXy0TMNDaj1fRArYX15f/pImuqgngX
H4O0KUXTjMPmz3U8hukre5MJXQ7XdIfaJyCPr6pMkL5Tl9GsIDeRWtWT/+HTb4E6rNGvlKXLRkoQ
uvA9C3NFP7WGX7lFc9srWcVi+QDdI0G35u/q9rww7GNL4Pe4Cp+sXFVKAIfDgtvvv6nmehXQhHq/
0swU4Ul806mi2rPb1k5/j3S+6805fFdofOwuHpyxabF9ZwbCrV9nXIi9XMUx+NaO2ikIM1pw1h/s
1lvxDJiVM2B3oYqjYHvwgTDdJI/Ww9FsMOkFd3wctxxp36cdGv/rpI2qGJVGfjIfjeFKlQ5NwaeI
IlNv9toLO0wdGQBF0sg3r6XQtfsQxxs6mOmjlIekVyQWQKL2+6/09obwcyX57fqLCn5D04dG2sMS
ZJkj7ngZibSv2ltQcuxDRIAC9beVBwPH8Az8uKZtxreJaYsc2ar/0haw4jNMtBkey+TqZXpqeCAJ
Vvaa3uSqBa0Q1YCVzjh2bpoIlw8lDJsqbmaDR9unqU289TwNuKRKvUiwmU4eSqp1B6VdGYlJJY85
yYcMIHd8hUF781/ZNYAoITwEFUCCiV1Ysgis2udCnzxpXTqTx5j/+1NgmxuwR+WFWsGmTXJZCTAf
EPBGnVFIeCKwP9X01tPip+5XMjdGfyuB6uVsDtGNOBMVQ4SVd7DuxUdv3yeFOV/jF04f11drFOvv
/m2iuiJhfcIJNHgnH6L2M9cEUGWYC0u7gA+sV2VTyXn4Vjbhoe9kaGL2e/UPvginBlsPbVBEFJ3N
7EDNoLE9iYojGr9CisY0tf61Slnecd++L7xlbnpkk+ySWgUlWqU+70JzHMJAnLfGIpmUK+sVzGoU
5vYobtyIEqv7UhO71jx+27oKN06yIj3LsZ8aF72ymjJl4utcQEp/ptrpWjQ/FC3rL12oC+iigfuO
+iyjQb05hpu85XOcELS9eMjhrcOSGnhpGk7pe3eNalfBej3A3qssk8sYMMKP9bteSswjVAVc4l0K
2lOqMvRPh9NQvNAj/d0ilurNxrWfdrtaRGJt4OIPhD9LJ47giTPOZdZ+WTGfduSn6wshB/Tfx7WA
TdR1qPbXMysYMJh43rRnI04km7fC5qUEMw9DzT/dXMJUtivfB+uBdEiSBUK4RNorXBQlw3W8KAcB
FUVcf3ZMHLqXTQZpvBYtrak7oJxl27+KJFA036yAewNhhf6OvP+3raILFBdXUBX9/wQ6Ty+tAblX
+VpzvG7fjcTvtJ3HVHy/fUbtmeICUHdcmlusfltw0tuLIukELaiHmqWAGUoRxmNz15Wvo98CAmCE
HeSEuIN+Kh6fnwSpzJi8aNiIvb3jlZDb4JpBKhzh2M+QyKfyyy11eYE6r+t8G7drJuLvNk5PLPk9
a0atwhLhkLr1fxmeGBNjXesXtGP3bBaLqyOFvpyddgBFe4DIc8ipHtu3N/jHCbpKSf7ngmaNRNav
CkhHUKNyG44l3Q0jQ7rCA5RWUSCdNfVuuoinf79vIDUQr2CyuBjLgeRhlyQt4BIpIzn4pSmyXOmf
qh4j6DTtfU1N3iGH4qe54W1YYsHSfN/Nbmwf2o3mUt/6BVycecfTxPmx2rKATfYaM7TZ1rqAQ7vL
YvFaIDGgyju07pezPf9kJaHa5kcJDlYgfv5mGrUJCAv60nUMKPl2ptq7S7tII8MJzt+Q6t0xFIIT
mWVJXc537UJy32fYaNz8bCwmRi/TYsxK+Zlf/mB/FTr4tGb627znOxyS+SmEPqmZrWCmGMW8DgMf
SZ7CBBipIBdgyo6yvMB4K5dwGYy3SduuDKUaL451UOcIS6LYsYuBn59JDB/AJ4bv+lr8Enoz2P0p
fmc8fbfwUSULLRNj8S/tIAPB5+SRe69EGy5jk9j+y8BBZOcL82lCurHKsgB2KK/zn7o6xHbP/JWZ
rqyiT6wIXTJaQul0aiHcWZHCxzYGNWAWz6Kh/sp+CkrO2E4aETtIGIHHhZnbjrn1UW18pacBRraB
2sfHsd641Zm4wf4mNMF2PYfgLJLNwrFBx/6KDP/A+hYItKXIjJXQlNAc7cdXO7jZ6uMc/OES9wPK
W4sAhauyqMfrKdlOKVkzNYUCNL/bq06zSLOm7YffU4+a+81dGd0d7o2zWR5vYEaXK8zooScphVox
xP69bzSTGA2KLrdx2J7cBFAxnn7SCK1TyNNRbTenFkpMR48XzlYMK8QoN8e7S2TcVl04DTUqk/1M
g8oj8k7O8KKCorqRMrjAN61330piBGkjKWhjUEujgbJkXsih88DDTN6OAwfhV8IwdxdJvXawVd4o
qDtbB59RHGJDnX5VHb2fsZCxC+sZYzM1OpcOr6IPIIN11OKEHgDBm9z41Q4cVSTKI53GdEhCdoLj
nGUy3BkUHfmdBBirpxLBePWmfAtAwcyUUkttSo0CzVXZHcaXiVR2x6E5PVmwnF6zqwwTP9hJzhCv
7iGdzxjFMHUc5e6aUGUUPQGB8alZFEImqjgn59h8pbvfQIcKdVaksGjvoezv8iMIQM/FvIxIuRss
SxP/EPVcnhrZU2AHDEnFKqVFYN0g9mGNDba19Roj/3OQCN6r5qKpgaMM3wlIYME2oMo8N9KKWBAS
uuWbdypFMX+9b+dz08Q4eF1At9qNctx9MCKAl9ONrnExp2FG7G3edz35C+C0H6NmBntD1HCZBfaB
VQL6EqHRwxwI4tHjVs00dmu0tSROUEKik53C83O0dbtfkwXebFludCKQ+CrSp6X2mbJR3Zu+y4K8
VaeDjdUBYTIZ5Ia4+Il1d3QoZ2rek1n8v3gfhMnUneJgBFMZ192cTUNcqr0cXp1JlAMZGJAuqKHi
f0LiHMzwSTrOqk5EMYKTCxk3PeU772ZSXDH4UwX4qkjiT4BK8M+r+1GVMTk5byNKBG3k7+KlDCj0
CuAyR3Rzo4ZraO1LdL8nEqQSipsAf9UtL/MMCgZN1pjTRkhyywqdYt2phriL8BY9MsvOyVqWz9L9
bcDDzHKiyLGP08QEAySPTeQoO4qWe5ruFz8KTWnXTXqgPj4ht+0Tyx3E5X168VpyusjdwclWprs9
05LSBdbqL6VMEMoZy2r6mH89KlZLJLoGC1JyDJQ//tsvWKAw+cuD4nooMFBeaj9hGNwQ1dRX6IVr
ptvvTKAp0GROM4+THp5Tm3KzmzXwntcORw82VNMHOGOGinN1Un5vJbbt3UDe/BZgqZ9JBvBWDAiP
Yz1xWkGi2bdP2UjUaf0yM/xJ9So5VN6gb2BcdoX1URnj2MovHZHmW0OMTLf97RynIK2BQl51KR6l
FX3t7TIu0qwyvCFET45XR+gNyjxJTiXrznvL3kR3bAlHwjbtD8unChXzgXNIcLGNf5fOYyrSqxX3
yxipKYYuLKuCy1qrPdKhfpOvp35hUFVVkS4AFX2s2aP+KJ/L7rzDQJ1jTF/DGnRjUWzkKr5V7a5f
zvhLnwJPJAcCUlDQPHxyiGi/RO6Zm+dOCGqAI3+2fTAoD8s4GAp+CmK3Ak2uTWadONRJM9u0o4CV
rKcuzMLF/i/Xdul30TE0MsTgvYvGSt6krvImzUHIh1597XV8yIld05njSWCaduMKaFZvfTXHPVPk
4ucKIqd3Nc7aNykdv67V7AW7ELSRGciA8V6NdTuYM/0d30I3tQz4tjk1k8l0uCc3x/Fjpan4VCoM
/iYA2O7HztS8y91uDvKEV8pydG6K5v67iTg9bnolLLZKA9mhk6fMsrB64EgVFF06h403rznFFeoY
pIVnRF1gVLNULFViw8x7v6Aj43MeEO456avObF0klRXEZiI0z8E67grRIpY9XpU902ERDPaKiYYn
6b645rlyYZ/39dmjJgwjXQ8rJ7HF+zIzuT8gM0CzyqZ1XGfBvKM8ZGpGuHmRa4KF0XLW5teIHliR
wwvUDnoCu70BYHP4l9BcMbxRA21+/0n995zqPkMO/CL9rYwBtSvAL4VyPJ0oQNNrNF12K34kxzGS
uMKQ0PzA2u3dA/QocqcEduUKv58ZURb9aZ5NtzBfMa1/cguJrkmmepawW19lRV6N5KukKhVVFFtV
5oThNV5Y7RxJ/0KBuetjEFhcF2iZn11ZwJID3pynyiM8KGWFydxSoWDICeAMHvHlzBrWHfXh60sv
ZybRd9ExvHfBfH2OpOQQ4jzSIRjF3abpX/QJ4/LIXKjjMdRFOH+yApeZUY1WzQ4By4xdgXXbqySS
1+fBsTzJ8XLffvbu5E9c4+CALzPVMWy97rDcBJVhjSFgEoVWHotNuNl5+e6FBS1ZBbSCxrnxuxUq
ALi0B5SAKml1odBuvkyHcYQIOFWaPqrJGjlYPaUtVxqgLLEgax/U63IlnG8yO7DYwQwMM02GT/ZQ
Pg1hb4k+5NsWdmr8BKP5Z+WVVOqTXyTTJCDR5SiuWTXQfZivABRIhA6JoByf2Luk/p2RdN6jtGZe
h7Q/w9vqLnCmwdBaoRbKkjQNN14sn3NTPCaQzDsAXUq1pAaxTyVZnLphnJ+XzhEuzqvc8Z9UOhIq
bt8T7gnFVs/4SUcv6KVq2d7SD1g1FCGetdp1PGB6QIsBdIlBVwoojxt5Ff2SXzPLEjaqgSMLz8Xz
GJjKZu0WAjTkYTM3bMptA09PJYoqigTIXzBZgyVDhw7idHhaNm/XA6OHSe9Q+w6szFaZFsQ5rpBT
aFlvZ+y+qSDNNTtAO4VATDxg8jbdbcm1hC8nOvpOzH2ROcRaW/w4Q9y4mTxw16P2Tf0KaAXbzHuw
8qbacugkwU8XS9eQBIEEHM9Hop+FeskJEFTt59HcKyvwvCOsVMXLl06zrGkCrzxzcGWPLxtEVGHZ
DvcIGECo7t9J/lhWk36RlM+UAFKEM8mbD9F4Ahd3ET+WWikwMKhkBBvKyiedFCi5Ppj45rwAJ19X
B6atXl7yef9S+45PIhVQ8LsRZET0BOCkKgH4+7jSGjrtIAlGi/4Xnj8HctA0YPIT1QN5zH+WZ6xT
X1zWiZxuNUYpFZOOdkg55aqRyI3mKtKHFeSt49POZOGtDxT0xKDTtd5mPz0/8P3BPoMS2UZQQkvh
yDChswyvH0/5nsC3dhV6s4u1wY2JJX0hRXSpBoN5iLhmcXH8KCXssvwWYIP02QEkoKIcExS0noja
lI8VHSZi8ecRGjTnP3C8peoAhA4U7fr3QgMHom7NhZzNS2nOklKyx6AZcSAnZC1kpuFjn62OknUd
QGg7WluZ26bAyn07336c5h4d+auw26f2KLE2X3UsC0ls2c8kUn6mIS5hjMCX3nrpmL/0uuVrjA1v
W23ehePiZ01FebpR+gVqGWv5Lamwz3pqsg+pCS2iNiMMQxnl86NvcH/+vbu8di/nUwDlhLo+AcSe
IaKPHdJp2N93ITuh0LgcQAIUPJXdaxNIG/vDJbs7fvrAGBoIs354XNv04YUTfekvsl6oqlJ8ukA+
0Vrq9/EjnObBGSWYhOVOomLnu8iC1iLfjgEz1VerIjE4FK2wSsN4cF6iKukylc2mB3mM1pIrkKpc
phJYslCUS9UjPQot2S+Lm0HpL+ay+rsJZmOsFK54CxSQx30jWA1amuysxr21So9U3JLYPEklXWx6
xrwEjgqrEcZIQFDu9ncFBKfEZp4sSMCowAB3KCeEy3x9Tgrpte8D5XMDYJZA3cYUz85hNEBGsEC1
hgYq0+yJDcG/XJeqgtunTZyrgv2E3AAE28s0rtHfZwXDgROHjA2nlIs8sv73o5h2HDMoM8hb8pxD
BvMB+CruYNm1StR8LzUruKAMcreaMklB0I424DcobKbjJbDhFEQu0FF3EBE93TnEX8Xqwlm1hk2X
HIrOlH+pmb3ceO8zQkJr2r3OchxIVaXyneg3JWo6dTIN/m5EtzPA5Z3Lw6FJZ3F1DrVx1Xgdla1h
v+C0L7yObiI0j8B81n25UwMySMf2FAv/Sni4Z50s2rGJa3tBBfU0+o8lEa4utE8Adpdd9wF3zxql
ty/kEFOP1c/w1cpasQToHuZKSB27Tg2cCrSwEA4gysZoN3Ht8H+oFbM2KfY8GlqIJAXgeP1B4Lua
+bqBzATkrxLH5M9j+BR5J/QZXMsV5KgdxZo8af71/ZWsL3tIpmiTpUofTtE9CI+ByaD1Uc2YJ3eE
KzU/b4LajXSgvjkEDhPbGRqeOghVmloEEswEjgcsEOINZ3SDFFNueFqBRjkyvsVlWxV8isTNjH3A
263L91cCGTj0yZZcSBRKcez+3s2kcYw63G3u1W/GvhvO0ZVeIAVA5S91MuBdp8JoRGmHECOMVcAB
8dHnClntN3yCQWeCyFb/e0ZztBjr97SDLCvSKbJszn3rT9q+rVXwxDUp/rUnmKvc6gk/ddueaTKf
hovuIB6AOgQz/s2jFNdBCqiMr7JuOEXdgWEcAF43b3RCwHuMHkwqWlwrUFfk8xF57BjDMb/3KETx
E5pK7doO42qBS94NVuLBFHd1gk8xDOPWar7yTE3/2wZJFwGDM4xmE18i4gKJSvsHLOgUFumfL+1m
sO9LDruWonFNqLNKxkvVUflOeq5SHJG8vH9HAlEbUsp/C6wUIUUboChvgkkakP+UUwgBOJ9DPPMz
6mfCGXhdBCbqYh754/gEz8NlhOaBytxzDWh1zYv6W7vIVHwM6KUAI/kkSYGStkFp6HUSh3uNaxd1
uzt+8bEmyR5DqaQRq9QIdTe/h0yDRvuK4iWGetBPOJ234zE1onHcpc6okU7ZHoCTE8LZ7zGz6vSM
coE+x+MrTr43J51bYT0U8mb1XLnZaUcQMFc+Pb24o9m5uFSYpoNu4LKmqxvnTQf8pQ+bPPvQEKF4
QnPnzDYMTErPWM7JWJ1KLYbEMa4t3y4Ffbt2P91l4cydgDTvf/sMTv7d8xTBEbntnSIdW/yJnjc+
Eal2Fpq43eCZgGeqnbyDJ9Js9y/oR0jV9kOSC2sSBJuDHv0Y3zVoS8/szGIDg9Ec+AfFu9CF9gQX
Qglz29Ra3RPe+Nj8mksC/VXKjzQWTBegwvoJor9ct744ikGk52zMAXd5+WyBbqx792uCBwmbbXaP
6Hb4AjNTH9eNoN/kqBXwhCmLY5BqRcggnZB19tFqRfaQC2DHshnHXcBRzVVbWaDedM1kf1EnkGC0
UBfsG8fvta9TYJVBCxDylyBQuFwJtsQ/YfOyoneWD8/Sxt55YzZQWRAHUngRILb0C9tBiGTxmNUm
qTA5erKnmslYYUidePPn5Uop5kRp6/0Gdn4KRrE81BqD5FtZFcGHrNqSLKLmtS/aknCh+n94+5y3
EcqS7ySqfASx04r1e8ksLNhqH4+S4jDcT/i7iffaOMVDr5k3rnnlZXRr3R+ehzJ5i2K4Uw/F3vS9
SfH9sLht+6WgLAkUqRXTiBaqcJBKS3rr09K5K7i5256htFQ1MuZ3JtJiO31JTWC9GRU+XDLFoCQs
cCWTn0mVXWboqPToW0BR01l9BK6+COMEVpxIxFXaCgaJ3ipbMnyycsWmKmNO7UN9MqYjFI1BKiCE
9y09HE0YCWymqReHDJwOZf7u0X7LIq8RLZa+dw7rlLKrmvDzbG+CyENrlM5bichAxrGrsWqtjC7V
FVawqut+D1YCXTqKbYWMTkPj7SnZUlvubyunwgFbYHt3Wpo19HYvyXrtq+pZeLp/UfXfdlCy8IWj
k9HO2SvvCJuIsiUBHQi4nUeZ6P4M1TQI/M1mxrAdyU3PnIreebAw/2QkrOv/AlAc2/9V9yow1d1h
Is1X90Uw4X+KT6XMF4QunFvJQLALgEh9a6wlXeyakE+W9+f9IVoipL8h1txznBAbFhFbshU4JYyr
fwwYwb9dD5mCGfS5OlrwMHF8nvxVdbaVP6DoJCR+25flB8t7irpb1CxFteBwXvKYEFA6rf3gklmj
xD/YqqX7HNXgt7oCy3dcPitdYF//bNBohwk7vdQZMbVV/8zcgoT9lBtVLluA26U6r0WQQoQWyHVR
ONZzMHPvBPoJDEV1sEOdLePuDD0dqeXN8sQlW/ilc/rsmSZgFTxzPQwK+x93XmeIvHPcaVAgChLw
ANqv53IVreTYDQh5jh4VnW5z7Dec60oocAZZtq//9RPkHhpkoYGlqus5GWaVoN1k4XsliKLBdAkh
TtKLgwGAvHGApv1baP5oh8ANO89ohcnUo0VExY6Im5q86KFtWnbuSGVnvGGu1VokV2dYNhENKcYe
cYSMf6hGjmTdw8jBAHu0zBb8xYYHlANrm5FI1l/iTxcBbDMSBSM0FsgmDSwUKn5pEXim9BVMIm+i
XpsYUN4hbVKcHP1eh3cBVnD0U+0q2WmWVmmC9Eq3x7KY3cDvj+lfAEnq5P/E6J7/4OeU1es0WP6t
QVwXzIxvlCc0yo7Bf8bIQ/vOmEk66aGVsFey3KkcWKoDyYALVqmMEqBendda/CsuZDts4HdSuYe/
3jU5zwwkg0HRQ7xLqezewDoP2LswRjVJ4ov62WGVS3XI6JFO1sYA8dt2xjVfy4LvnGKOHHr5rADj
ByuAO5h3v29e7lX777YXA0c6gHlxic6o2v30kTe2MTUgnHWJGFV2FUr5LB9gc3DNtvV2xrxEjPNV
HqoeisTmnSkJZpSeZMn/bC4z0zb8XnfGgZ5xzP9CWJW38hu7rUhVCKLb194O44ZJwWirDlRx3dHu
ZbdIv5VvSPcq740dtlxgUg26A1O9IfjKmrfggpesfHyufRe+I7AEhR2ahpntVnLD8DLAxksjxYqH
Ca4Ff+A6tAUqG5H56dQRE6b7jOvtqqDm3kMy7XwKng1a36pEmJXnF1Ka0hJJIKp2w1rn/ISXUAoV
P1N3QJGEd/qWoIs0FdqvIhU1OTBOhskI2jWpOYM76iLsX2lqe9D6NASiR4WqJS+g+rEUiyhJNjnm
Y2tqe2ySJCPy2LO7gnE8R8ZEBMOGtL1mtOluR7Q9lxO6LVoX8WjHPbEVl8lETysT3jl3dWg9kKLC
Nvxq/JhCu9g8db3LXeq+SXxC/jKazYGR8crQPVmvpSmoqYJSu9nI4Qa4sDEpGCo2RwZBqwaGbgfx
h7i0xvNQW6b1s1/udiMyq0eJNtPWwGu9y0UY0j+mOiG7Y0mY+XgcI2grD1vAsBNhUXcVdAKAOs0K
OAD3CSw5CfGjUy4V+69F3SPMkKADUPn7KNByr9KYc4gHaTZE6Vt9e9OwpWqFM3qDtXprGK5k5VQ4
k4Y7jtLY2ukChkzKKqf162gh940cXC0DbLlJcUqDSPds5GpnkByrCp7UutQ26fYuXABQ9vwkQRsX
e71zpv3T+iYGL97zWiQrL2/tLun0jLow276hyAosQCukYZsVBcdbEIo+Qub9N8npMhtXaCs4B3Yj
bRu/ub/KMEm2Zfm9oVd7acPx+KMyGXHLgDU3IqInbxKZF9u3zVuvMyj/eDam+AnHcI1zhVWwZbVx
G9BqX8+AvEkNy/QqfJ3uA5o2hLNnJqMI0BwJj1VaPHVRElPCUvl87mw2LTqLWS/oaCx5wxy1JZcp
6XNI15YXoRNPn2O96sxjmeds2dp7rk5cXbOKhgkNUlw6Vd2CwYetGn4QFjt2qEP9NzNQzMpuaSL3
u6yQmGl0t7NrT2ZEiGZeAnRU9kOzbKjMIpK7LQUNaFTHhqQSo876n0A2Jh6zO1Kda3qdjvrqNJUL
OHS6ifADn/Phm0KKVRzlDsGvYKYnAhz1qe5deQvf+b61CD0F3NpV8lvJY3Mb9zGuu4seCiKrrowv
0Lk2XN/Pdg+KHmq9dTeKJ+bw8S5qk/DXWR92Q/9F4cpxtucM/BhzTiAovIedR04bU6en7C0kzCCH
JSsgY0Yb2ihMKSxgFYpIXDe83BVpmSM4GeFcu4oRFIVqEf1jJgpLripPaU6Py798aTezT4lb+Yx9
/8vj0orr6paYEg0Igq6znK/DSNNWsvwVE8jSe3FIiGw40nACwgTgCo00QVRpRS57+9ixR37uMkzK
++RzeJYZhHxlKxpgpqC1eWTOw9eQvpbSY9t6CHNo/piE8g25IgHW8YbzU06g1se2PsskrMKN1kut
+zewGukXSCocNEx1BlgAM8G/qnDlSxzwNGebU3U8xMNjx4440cU00ftjox3atNBrs1LI/UjcWidE
8ZFzmK28YSnW8OL5LdtxO23hg1thl8KwnrjlmEf24BskDIsHr4fkOHKOo/eyc0/SGLGAa5Q41WeM
c9g75h3eiVkXXcbLvbNFDfxgOPP4PNciBLJcrysqEstPMHEjLcpytnY3nqAQwAREm3dAgimuhL6n
QM1uPoaEMWiF3NOds+gObP+YgZxJ1Hofmw+Z03vFpd4lfeH6OpfhhEFMJUDT/dTHKIYlwx6BedUe
lBjLXUa5CW4OAksZ5J9k9TopO3jOdvOTZU7JR4MY3inTP9Vt5/4EkR1lmZJlZF1wmlptMDN2X0yu
bSryFWh5FlXHkZuzMsqbik47VqWXSrxe1CYfs36blppPmp7F1C1WC8EEh3YIELchj3Jj7IMbTlgD
5g3OuvyyZ2Bo9fQl0rTLWjvb2d2pbh1DAUcrJgHzzEp2+HkyaxQyAOi0dX/zrCyhF4+UtaD0tmxq
e57HAvhn46QInBm5+9BcGZL83xqC6XWJLlJaj1HLZcw5nDoQlS8ua+CROJyM9IDyMQldVrQLHbHI
KCU31GHrl+WGoC2NmKaceOgrE3uSTfmlY/SyQIbiXc1JyCmqem60ZYJXAk9wMnUao32Hw2ZRcAv0
huujIs14O9qAfLQyQYhNFRrOgsURWCcR2ThJ1b5WnQdquIZkvWQ6aYRG9Mwy57h6Jicop1dXD+Qd
+/YbD2LnPU0Lf3yv3HFFcvseGKzL6bv2SEadIrhAv2UpdT43sieV7KDqLmiVrghO3FXMwU09nL6Y
lx9H/CHsD/DNU28aRBVc/krnOOquBdz5ouq3xIygCHyBCeOc9wiPhftT3WCCkzViP42QNPXj/tzr
ReygfJfBnwZ6kAA7oFa23mqUJU0yGLCuHP51cyQmo3y/VrmM6kT+rg1XIdOgUIZnqBADGWCh++S6
K10rayIILxdGyP1WnFAZjlTndKWC/yz7E5yqUKiI45gQnXxowqHSnZT/RRIyBdDiHP5c52f7KYsN
a3ujwZNhQOUQlddv3pNcWFWlX6uh/6GzrZXnfRsNrNVaG+sd6AeyeffWR5FSJYTSELHYdMxBe9uQ
qFchuPRNHDtMRBaqgzUQXBR6Uy2Z6m8Se7xQWbYfMMVqhwDXnt1tEvVfrbuiTEm5bqM4+jfW0h5u
phqlS3xwugxqC9ueFyG5v8z7O1UeuciwIEXi2MzZ4du+/IWCoqB9+pjC5VtFQKUSYX0s0s/EtwEO
/rv56dV/eTnWFmkiZcitCDVzk0RPGTiKEa8x5pOk207+acqcew4ooI8aRXNhT+AjbaRhv+LhskhT
Gi2xHiG8dUqSdM8=
`protect end_protected
