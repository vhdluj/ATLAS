`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
X363KK/wDFDgUICPflqGIkvHjP2K0rliT4wb6peQVDwwp1GaSKyAQlfusmI7gmDki97j3do8nwXi
y3tCB7vhzQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P9GHhthJFXnoRGakgsKI8j9tgWRVI2zzuZ9D3mMF6Y50os16HHReHkIHtwmPn4KVSdMTIsI6J3LR
gFReEj8UNze5AjqkwRKYpDjExcnSqXAmcK/4M9u2gMji8zwpRpBSRrCvzNGYqvsXFhRESjSyoMJv
RS7RtxqmyIs1CTDVDMY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t0fXMJRiXvhdnsGGDonWmWGRRQ7MQXW8xDLEnE+vm/lryKlLwfqXEa0vRRug297ceQ1fhOMQvpqA
cLkHTmoFRQppgvUV5uDdlhbj2sQOLT7ydbgwvcmr2TzkJSZccZ1FBK5i5cm0dURQmJ28UwmOqAU/
nvbpNCco0sUG6sQoCpITw4mH5dRk0W7pwpO9BsWwpTEb32jK3dXnV+40wa6Dg6EPvS0/9WWv6aNO
AkYcWnn1uhat1Yp2auXE9E1A6Fxq1LOQAfDyxR0jn25p22FfCkqqmNAE2aiD1UYssXZu2+Y3eurh
UHfAs7mtoKXUq/5X/b8AtoIomxp4Rqab9ThN2w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
npDrda/gBwvby0iGtOAAwEL+TEbgRZIpBzWdBgFgHC03N1xyJV6UFlQC9JjKXspJ7KuYyw+hxvyV
Ap6QzaOT4hv8FTTutTjvxkh0fArNdcz2n1VOVq5QNnmkrJ9WW1rNcVXBxoXuVo1J03Vh00r/ESQ3
ICcPX89q0+fY4cUHlEc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nP3qGb7qFszh5iA8YQQ1FoACDElTKnawh6W3nsgruVUkRdlzIu2Hkt2djPnziUIPK4YyvbLMx/CU
ux/n9odR2X5QlbA/c5QcBkkUiMK+87kmiZd3wEdnj+vyDiZg6W4ghEhURs6p/nQp87xM5w5L3CP9
UPatsi39ZZwaWg2BZOfYSFDMOLRrR8TD+zJPv0WpPHj7wwL722s0TT9pcKsHQxpXSPjTI+5Oa/Zx
+wGyfq/lG8QL/r3WtiNPf4Cs7APVVfJpz6040G59uPafNDNPNhKciuCsixHB0cthfnE7+smtf9LC
xQdlxItc75I1rMS8zXdmwZVMZhZLm8hhxjVv0g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24496)
`protect data_block
XVTsJDaVfaMxAGaTgVakLN47aBuvDXJQqdbfoy37+u/CVm3lEVpwrCqT6jVcRqmOOctwc6oTP2my
Q/IW0W3WAjkYQ/CYjI0BRTGvHeXIFiW0XdCqComp3J8UrSeMnZJCJVpPM027rVSFmRp55X8JBw/o
baANWnvEmHkF87szH9jJpIeGwJPDYfmb2FlZJ9JEnu8N2iyDaQARZS9FBWYIUlOJlqNPo4J5TeIk
a/U5yfZ7voptkkj2NCeZtAnB6S31yAZkWZA416Zm5nRdNHU+VaHvszOzDWPlAHwTLwldj4RWPVXp
G4lKgAKcA5Xser1OQdbfByUdZAMxzEcwWlCu+jWsNi1zFqMlu8j82Dy3sG4jCWeOGaM1Ex8WcMu5
1FSItfZEvN/pdwCCKyREZdqIRC8LcSAj0oOi09TmfcGleur5cfO5ZBd7PUEon/sVMDlkMuiYhNHK
fkC9pBoegs/2bOA2IrmowL4YAOnZYH3KFA1Oib+Mpn2lGZwNPDGk5wtZ2GaW9lsaDa+qI3ubsAuO
o/DagSNcxDPy8MObk4lrsKbwodZjsRO/TF8QaVd05Cg3Bu0sNCVcX4nGlDhFDMSbTOHFwjqL0MfA
+CrZeoCJbwMkguH4WqHzVZ5sQVXHuGy6eHWmLgumVDhcV9GiZXfBCatpBfwEkLPNMqIq3LcD6dZD
APzTXQZlcAvbqn6l0UZ5UVnSP0zlMA0qL3cRHZBKnw+seRg+gub/vlq/dlpkOlldxY5aQmEg7MbF
OOK01Ye1KjAUaiCLNoLGfSRgmmOyHjz0hYpf1CRA5qo3/vew/T/wEfUWL8lnf44uRcprNltJsob5
PoLIM3iN+kqHS0zz9XhCoAZo2iWChEzTCsLTnu9DTT8iLIxslFtSxiY+kLKDJ4+NYB3n22yn4+9F
fi5SLaMajqNxeoMgtI6BskE/MQ5NbAlYq8GUSvi5oEx3DZ7iYyOmiRGueLGnNmCxZRELbKBRz1xT
gBkUvDXh9b6Vl3jAkVzqpy4jsNG2PUg8I5ON4W09QlCxLVkirW3PPWja6rBeQk4aiH6z2Rmd4xT8
KT/6KN+S4TV/iHbmF5rlOISmJb2R19rIxENO9N3dHUQLkXbQIQvyAIS5e6xaG7pBRoW4crA13X8P
FPO3Dwlr5RDrt2WfN1YDCjjUinUlfV0WLtCjR5X9KBniNAjmBq0i52zKgbdKb//ukbZfOjL1ereE
dv3t4tHPOMwcxCvSeL9CqmHCFitEoVsSwQm26qPrQ0NxKQP9Yed5FGP/v5Z44ys6d0ZX8JJjXUSn
NGQNKpb7hRNnNXocsQGZalLqs29uvMRyydVIVZhfL8F2cL5Bl11ERNbP5JWQczbTznRDQYGItsKF
Buda/phI5MzFxkEUwGH/OZbpgckFIGW6r/DmJT9NLoaAB7Rl273ZjD30vXoQCMZcjYjoVnSvxjA5
YeC2jQeA3P8rFzeHawmDmOnTN/6Gb958dT8c4+SisVIR4aCmyK6POtj0LhjpfTrsmL7NJ/KHCbWX
Ai8/Csja7W85JxKXe/t5V5wP3wac/obWCSKIjDBtB6EtcaFx5uEd98XDVSEiJeFHXkF6TJNKUesL
+IeX9c0IgIgU8auza91zDCCTvIwXEjgecWPldDWHfrZ7voSYn9XYUBKFyIIl5/Rwq3IamfUNcCh6
gA5VkCxkOgPO9JgG8jmS3zx/LdWAhxEntQqnid8g5rrVHvoNaHDzCpWQHbh3sy0pKM3P9CrIqoA4
41Gc/VjObA4MpXz+ZgDAvdUhuB9TVjxczkz3eiWHUhO4Fn0R40MbJaXVM5cabemYe5FAw/s9e/51
3jMpX4nW0v9+6Wl5pG8m32fsI0hzSb/nw+ru3q/UAmQuciMb60s6qzAVV5B4y6GCIMcQ0by+7yNo
mB3OelaQXY2VMSimN13wuEmhi5phVGk/g/UXpzdeHcmG/yej1Y5s4ePSJsOEOpMQiR8Vhbd9xrhk
ImYQYv4iacobhFcmG7cL1CjCOTRQTWYjFvbCR74BsqOevjoY4x2N/NGxSz2ZetGqkeEEprxzD2Wg
4paDzLYdZqeEOfiNScVQHWhpipnbd0tsUXGpgh6BiltbJ/p9gjTL0dsmLYzDr2YwtcyHcJ0cCfM6
U6iksO51cREWalYeTTngbUE6/PrA26em1AMwUhPCd+guE5wQTOtOepo3mFguGlbAe/Q98kdIJtGq
WWxus4Sk2N13GQ/cdwHrwy1zWBy6rpe+7XGpEgW5AIvFXCoUsED7VzRhWscIitTdlDAz2lOWm6Fk
/6vLt2BH0iflSkF1qjfb44+FkbkTiahBw445oexV00RO7SxLjeGMXXGbq+DrO8sNrHm6Qf2YLPDg
fY6wGWcvbEP7EhzCu4lB4ddaeCuazWKm6YkHR+TGFJsN44CxLjMsu9x7QhsiKeQWg9gxArZW9jnY
VNzmPx8zNwmJmOEpHkZdvAvxlnNM3b+n4qBFBnnqyJJepG8P8A/gLY9zuVJOeoF5ZQ+gDo43IifG
NtjgFwuYB20szJApeKUhotnCHvW2KXbKnMxYj15Iuj/Wx8bfC3bA4TH3Dxae/rv82vJTzBFObORw
MUN3ExvFLKIq3oX2RD3rIt6skwWxsSOvNw7DAJi0eoakpGvL6nkWIbUv2fTDkoOb5VwcsESk5M2d
FgIQHxBbTE+X3i6AtgOjuVACiE4AFyNbUFtIRrdrxsQkVZwhC2IpYPZoe3RNQMie03iiHCr0muAr
UzP1eoflHg99rgS24AlVWq1pW0wPnDLB+MoUgrpNv4oWFyscQ3F4KGpueHcQOw1bs36Y7zQAgMM7
iqo0Z/GXkrmzVVWLK0sygInqI9gC+YJ3iLMdlE6UHY44uCHtL2EG/SsquxuGNgcMd6N7fHmTKl5e
91CyZZshMXVdxiQP6XWx/17itD+dmaHXmgJ+XMZ/lU/oBuZbnukEJMlnG7q5CgKUR6aAvOV3fSTY
N4SdiiHfbbunT8ABFuDUnktBKKXgg+q2nD0OVjeHH8tJb0D4CYALZWe7IIy20le8BOn6VKv1krKE
9YpYavdf4wFrp+odzPJTeTnQY70G/yFNezwwIN22k3phEmfQH5MpT0cFwikceUkv/AbIKWwLUJtA
+cvlWOY0xL+Zixe7IPQJmucq5NivBXUYMyTzng3hJpZMYLWUYuVP577UtKSR7alC463K9RrmsqBH
tTx2r8qx23DDUL/vwZCo0L3VNi5c9E1A2uWzM/2c2lRUXQ0CX9Jk1Lx6MMbEgZ8YLgziiyIa153w
KfzwzJxIK9kx6OQxUeWA/IzXpFpah8aVactVr416gelS+nYoVsKFY2rUoXCbaKLmbgLNn7Rdyj/4
PXK8vufILPwOqoTTLMBZyq499S+mLq/DpMLFVdtGh0vDYsB/Fkz5TPYJi0TPOgFbjxmdRF5bXqMQ
hiAD5//JnUMtowo4CP7ZGisKZZ/woASoI860Q/khSuOu2E+vD5Ytvu6WHZZCqjGat1X6QU8igW47
KV5xOzDHlMaZsf7vWFadiU3QUz4wgD6YL525xkRlEE9Wiz7uJ3W0y87DpLWIMPCpZB1GHpGeEuxp
GME2Y2ce3VqMAa1QSwnqnrzEk30yUPRatP1pkNl3RgSHzHoAHdsVGie3K75rix6oPp//CLcfbMbk
Qkwz2G7snXw+uUD6BlyP72j8hAYmKjQ+Qlhzui6kzdCPphoutW+BVJFYX6xHmzoqtEU+Oi8d7R/q
jMCV7SBNVdOima+N5y1XeBpjULepU81drdZFI3qX3KNcMBbMNSuLyLoqYDHvlaR6/ZGgzT9yBvTO
eVw66Pkca9sUdgpLeCQZz9iZ8qzzxOS12fNbggv9RsPQr773rewN82lqJM/2ZOIPjes0+T9okhix
ane+QXPBsuE2eNmPG02VYl2CVKSvyVzrTpGSodbNun8E2/uS68olnDSSBbIqAqrS9xeZ857Dkz0i
pC06KWq0b5qutQp0ncKVR2OWub9smflRQHd89ZJfuyuStgWwopgEa9FM93mabWA1XaBHPBRrmlTO
eDQ/BJVteLG02Wts+USbix8rKKoe9LG7yYnFeqQht9k/pKvfSy02lj0pwiJzKcEEc3zdzHLanH7f
kmu/ZgrY1q32MNVbltWfopY9pKtmvxVriKXAmXxuarujbmdZq4P2ILCqiUqkWae2WPJ+ujN6Vnis
lDgiVoGbVyYs7/oLNBsqPcdodA6OjzAcdcU0WXVDurfkcZk7thRJxjUNn7H+P9/gCARMONj59wcA
xvMUoM5r3DdCN9uSBSTBtbs35SN0AlkUnDx9HBLBtA5kHrL5I2a+RmYTpcKeJ1j5HD6fL+fZIoW0
ZsQQX6bZu6EyWZfcEfRr0ptkLpda7VnEbghtgKeuplzMmJ52rmDEy89N6/V3zPKE931Nz8BH3qcA
JRGGhUuJI2B9wKjAJOO8mx4kdFvKTcTveD+qSIAmX9sKaZW0bVe+HP+mdYHTh0I/q//nnvuTkbyh
Ho8M0GKvAvZSUDEQJ+joZPexg7Ax7lhFDoJVh46Bacmqv7GiHxDbz3yJaXdiLR9EZUDQdicnBpCI
DFj5SWhJeNOV3FDKYDxbd5AxF2RqjZ9SZ900wTzJUSBTVJHqKadreeOnkqzqyTV2kwK7v3Vc1eR/
l3zuvU0ESfhm361AQChAS7+s+Hkq4EBRuNSRBCV+Sj1Wrmav2tajyBpB99MOEetXyzPU5TkqNjkQ
nztis8XZHHFpyapV9jLqdxHQWm7Z2/bngzkWKihuNabMOK+GbYNsH9LeY0U4pfvQNftoEmZIvH+M
yaZEqtbpkqpiJUOLF2J3TU/aTS5fLdjspi6pGR6qiyZCxG4qu1KGG7dsEh+LGQNHZtvBIfcXmJds
XVIzkQdd9n5UYHCJHvLXhXEcy7aO0l7EzWCoCzid2vtAh0c85VnmDpQEhheV47CYUeccafD6gD93
f4yfv8CInXgPhy4WznflixDxeUl9DG6slB2pB1Utgz5Kj4HIpsYBgIfIU09kCAA+A7WIw20u3ROs
8kHWLwleKnqmKxuDZMKCrV7jvD41bBqlstOUbRYm7RKkg2VN3WWqBeQNHZZoS/6sIpoGOSuwdWU8
HdVRllSSmdFCPxZERU4XIvh9PfVBfG1ImraVRY4aRWpPOTUUn0jBXsJVukJYRTOmOkDZ1e1RDX9Q
FHqwfmzGqg46bdk01myD8AE1Y8GZBxOMb3sRap1OlS5UWcQ+emgIQXqHTmpe38qJ+xIZonPS/UDh
Ob7tdEEpOk/LSgQH2hDGWKZe00dvnl+j7oge+QtRYQswfCYEgIQYmsH5qd3IvJTROPnvEFmBfpLZ
qg987MdBO+ZhEsnFrYr/NGGG+l2GqWhrrx4wuG6gO2q4tIQnj6KKgZn/fxeHsLoOg3dUwBN9Bex0
c3pwk3uzwwtMFtF1PziTwNRP5b54mSo8z7HoyqSGw0OPuqZPWvUEDeJbNNZVJYknKog0sYJwstna
0fM9KKYOLj0tVfqew53b1Svk5LfFAvo1pik+qprcPt5edqoz081xgWbFi4UtTUo4Jy5Gzu2w8fb3
B66VEy7pug9iQ4gr/5izdvLN603uXlFX3nFuUrz0roGs9FIF3YO5L6dgsdiYyOnXKT5eB298AyzW
t5e10JnJmxwW7wm8Y35+YyNiJr8mSmyKOk33qYA3glhlo7tXSKNBpnemZePL/ByK5DXWaYE3N3xg
3YAq3/VVcMlELQbXU6kKyV8ileDNWWc4nNiPTASo7SRWF2L601Y9ZM0trNsZiVFK6vDSOaKNRxzM
4NLtqbnYt9nY5Uc+NmJLNmHJnAACrlDtSPY6sRnWRyW8y6wtDjhKJpA/qADmP6Y/sgCBJDNzQQZm
jH6yrtgLAV/8ZuFg3ZdXnXaeQbuD/UwYDaFlyGa5CPXBxFEEstCftLdo0+qxBBcPTrdYT9K2rTX1
SKPUu22bBHlNY8rCny/4Qiqv7mczRnuxjpksOSoCJ/u8B3IKDP//UEaBAhOvoOfOj8eDsyW4+Ouc
ObYYpMhmbvn48ZUnihDvje2nbNEahCfDQwlFbS2qs3Zz6J+yXNx+zkRFO247LTNa6JSDK9vd1RPU
xWC32/X53PXpS676e/ozWCnPJCuYzwsAt5yKoVPqcM+XS4+Bl8xKDxiDHHu7Meg4otpPd7A5ZooK
3QAgNsQGsOdHmEEpHzHXP26wfeWLL59GTgQTr2dcanT6R+cvBnizSjyHh9NpAROLMWR8bqXgkptj
ohIO3MKn6ynUcBtuDtQy4tck8rHrbXq9pPUQzSNXOfLqytRPk88w2S6McQgo203m92ttSnEkgu3r
IKK+ZQ4u6BxacUKwtnDLksrcK/d1bAOZGepEk/YjgnPgTb0DG2IvH6Ulp5A8zXZ2bxrZxzuBJ9z2
7lDwsgVUSPYFo9kktXGpx/pjJ9a70p+fKExXBVKF0h2yM1WFewDJ6XoN0DKNyLFX2h6lovhanOEc
gPdf0YjtTD2gMmjYsgB0qX6mp29XclD2MothwBFKQ2nlIWCW06IKYNLcW67oVFkFxFjWsfaXIA+p
tqv5EGD2DW0vDzsapNhwVrQnEdIP03uYbqa4bFWAZ/24ypznijt4VtczoJwnnw4FW7k3ujXDB4kc
MIF1K8tySP818gitdH7os/ya39VFLbuOdfxMT6IekY6I87js8U7ODLld8zFbs1aoE5ztYKNR/SVM
7RNSE/V2rm3xHmpJCFtKclcSrcyur91Yv4Rqrnz+n6eKhcmZNok0Pxx8qeg5gJ055FkZhEcJ1ddf
AiINI4/3U5Qi80CNH7hNVLM7b9p9Byzx3h4Y9Ce46itVPB0tEq4lUJ5m7KL2RzuDPF4kJDjvHtcc
92bBB9U76Qq0qWhDMrzmJGrHpLKcvGhZF++BfPMELTjak20UMTeYWfNX7KGA52JM0WU8ZBXdHTqs
+aGmj0ErI9191MXTu4W8hYyWCKa02apHy6uRGvlS5E1kWKjDV4HYC3c914VOCZ05dN6zpPrQ7Hnw
oqC8kXUYkc/HjDzckuuvuN0fLZgvhVdweIyzraTnKbrRmqCaxderGb5O19ON+klBpOqwfM1bKNCR
Wgwwgz/nvUZe59x9A9vflI8Lr2d7/s3bgHcXZ9s7e2QRQDx20VkLPjFbgtf9XXWwjLGF0Kn629eY
wccMNpYKOfsdUerYefhIg7HwQ4BPx+oaWlZPCNc6dTXCGtHTLl0PLA4fYRxHSDIf5/+dGg0N6H0Y
3GLV2lZ6FCYC53MATb2Y+bbmBUF5A6L6Q+4tztORotIdkxJcmVf8aKWB/DpWQyMdKaaP0Ygv6ixp
J/Plqguc1qYjrdoP8eXB2XhgWoFU7gqxj1n0VsaSY8sH0XfCVa9+NU1LaW4gEac3W5ndjcDIJOt6
ACh4C5kb3Jtm1RdwlALaF0DD1HP0lQkvh+eJJZMxPtJP1mm76RFUXyz7O6+JiNMI0ae5rOg26x/9
BakXD7I3PlpAA7Ci6vusL7T+tvsn4oEkN7c4X5qc6iwp/l1dehJvZjtRTjYtKVThA+faTQLUg0rC
7PExgNQZ+RE+QTI0EKtT63bwXnOTY25kj/2lvRJ2bkRfatNXhh9ovJogbSUUWPFgA/+kpoRpt/Gw
ELJQ6VzQ3+CpBgTJfnZzDXy1uWG4FRyqiFuc0ROLBuLzPwWUwaqnv0ZpBHwxB+kaZ3MdWRabLD0K
qK0iXu8K4p8dCtYW+wtn/sHq7BWi8S5Bo/z+7nhqUO1udRP26UjebTdvjPK3xbJuCrGJ94KOv8vN
qXm/fQABB0p6OaKXRVM1SD3SHdcibdPAmHf1KOogQwYKsmyG5Lkk8oT4Qkn7F1OMZiQsDPLQ3Khl
JSlV94uB+l/fpUmdJrBD5U6UsVXnMmHB51YLJmEaGYZfUWV2CBGDcQnxNaDA8o9VCW/c3BaY5tAU
9IEIwnWHjDECl7mEWgGNKN4paTCy+DP3GrQJdNR44o0DSN+XeJvBrRv/VReAWUYfOd9c+rpA9+fA
TaO7H7745PjFN7oz4JeMCS8WwI9qLENdO5v6Z+9TP+az/OOewbs54w/gJ/1dMez3/kDG5zSVqFR3
PD/OLkoPk53BneU3O/5NpPBBdyhh4wncpiq4kC7oZMTNOInW9xyXcAbqJ5BUojdGEAzl/lwnyDx1
yvSsuBOiNavzOec22e7G076A4c04C0pdYbbdWCTzyskzgh7FyLqtljmWvSSEhRKliu7nRC72prK6
Ni0OX8c7k2VYx3jl9mU5XPKLa2tksf5VXNR6NWXgRkx/bqNSwMVmkqSJ6dSaPadqRlcp3NiGvYgO
SC5Cv7d6DPsGVPVFetkWWFnQHEB2Djn4LEYVMOjI7CmBMTm/JOqweb2IfuBmPLSlrYdnC2dTzifm
CDqFP/+8VHLBQkRsQyeDw4o9ZhYcTo0wBJ9pd7fjwiRBMAWGGMJ7bwnCJLxowRb9An9To/7vF6/3
tVL6YCTX7O9xpPQrHJdn1zMnJD5epyDzTqKVwHsEpkdCDYSh9msxD9ogcTeeOhKQlXkElXN5QnJp
zQfrJA0czQujaSPjfkCRnJ513NPcm02W9dGxpZUdjRNZLRMRSe6XOGoZC8FJvrfs2GKQUAPOO4h3
OnYnvaoWHfkf3mLd9UXC87z2UBGagtINtzwIuprdSuiUPcBwrd092eW+K+LlKqe9qX0lN223mYYb
eiUvZVg1jN2YuHciBOJA0ou28q+Q9I2uiMnIzQ1xMRIXlHsAGxwU4GT9VHCWKndCKrotmr5K9Pam
f6AQPQpOoIa4zc+/dDT5VGdo3j16JdK7mreEiLds1y3j8Uqs49j5azGFY+rqQNqiSN8uqDXJhzAj
5Hc7dTe8+7y9uil9/4yhhJnvWt70whRHY5rpA9knLrXKdYEgQqKjLdvzm4NiTSI4mu9XkK3j7rJe
EtwVKROd+hphNjUckM0PTaiPIjASU3fjlGE+FR33PCli5Wg9vXe5KyGefyOMMWDVZTJ5AR7xyczb
RuWztpk1/egvrBVtTbNNhCZbd/SRpjNArw+XRdVxxXFyCsCwJ512rqYcb2khIdxxps4tR+hVbu4s
MCi1rFnI6QynqNVTyKg9zoAT/qO2gs0762vY1ZByHb3QPTTrrvmkSiB/HjywTpQPZarXy+Ph2+f1
IfxOWZh+tmOkpwmN8Sqy2dwW3A9amNdz+lM3fODLf8lO8002/QRFo8Akx/9IcDz3h1GF7CDXBYI7
oF978/YDeXhzXCx+4iE/wKMWAFyQpmAMX2afDqcDSkQoiKRPgC6dlMHEfeU8NWGZMgEGhty6U6q5
fex0YhyfHu3uksFpypRAx6OnFr419AWPxfPCCLCdLWCJqe6qkYz+bhvzsLl8n3LfRguzyi+bLMqx
vYbDGcIrEinvU1L1xk2Q6Gl+ZSscNlsVW3dOB6c0RyfZhudZpsdcNAzxsZJwAoAR0VhcPyIvjVZP
lpko1KlorggT+z2SQ/uDhotNcJ6cY3OVTcjv6o0sWcEqPToonN7i1Afjmu0JraINYCbK+y9xPO7G
+hdG1C6gq1gHgKxWhPq3sXvt3Cu+lti/DZqLlL6lDD+vN5HNZVxkt1SMG81gvWUbItoBq2xTCOQE
J10fwh4ICeRIBt/4IWTGl6Tra2UgwmxStVAuWPCq5Uv2PGDfIyImXsAUrUKh12qJOT1WVvPCUKhP
L/wp1eu5JCP+KKscl16LZjCg8QaMWNbpdiuvzGlAnFxIDKRqknbyUmkB+u+KhX2gRWy7wouW1nsw
+XYhGTRfe0n5rSVH0Mv4P0VD6YVmG6fZd/tZctBs0Jl+BPLxPvzuydvL5UEQBY84VTAoIU+ND/3Y
I4X9MAd5hyuZal1ER7FaqyLC1Zz2TmD2l7ToTYV1hg2it9o0Pgs431T7JokbJ4S//YQ7UquV32E4
+/733hSY3rSn/AfwjPU30fdVDe3h/xLPqKVBXYiPjUKzJ91FmZlIZeSjntHUJqdbGiFAMKTjpdb+
zE1yvro3OnhRP+s35CQGnaBStjnuOS1N9W1AoLElmfGK+KeV9tAjDeGqndkby5NSPIYBEE6Z7mWY
rhD3cSOGFpA5SB8LBCDUpZvvsWCcSq9kTOpfmAhf+CWb3bz3deGSZKXemFYHqIHuK/FvjXXINkSf
qsR+di/WqdGJiSABbUKJIhAS4clnYy3m7ltAGHueExeIX8QOY/+MtAdsn+nf6kz/VGnJNnQvp5zl
85lmBc7rKVNaVnUJj3h0N1ATJoNZKCCAvP7MsrzrXyUmNKdfX0Vn9UVmKp95uQYcRS5Gjo02S0Qy
iSg8owMAS+BEd6GiLGSbEJSj7Yx7X5z55s+ngH45Ug/C62QWQybExXO8va89pjFo7W8BNqSQFsNQ
QOpSY5gfJqEB8qTLW83K1ULStTbmQxWHA6dARq+d9rwrPu4hyyx+SwIYAksoYXTIuyzQebMX0Q8c
vF0zKuPrvuOfmpbVFJ2hw5ceW392iShqMEVKqrO4EILt1TYSJJbSDyVkIXWMWPEUUg2xRti2Vaq8
Ht9YhVjZTwK4N3zHuMqnIdmbV61OqTMZTX8117ZaMpot7+vn/pjyNY4avmCyHEd+mp+40k8g8yuR
fteupTjNX/arg8a7fjmB9snEHO5lxMSVNl653ySuSJZapSnm9iJMVBsJRtQh1JxZEatjJMo49S42
fJ9YjttevdfmA5B0s0ipH2SuQZHWZJ+aFtIsfLPmaaAX706UjD4Hn0c9YMJ/046VxRhrtw53raTf
XPrPUSm0JvLyvuBcAhUKp5msZOmZDgd3Gj7e/uXV8twTUom9m+cQS9BKELa3kV5NkQB7j15vI74f
ssUX8X2mZ5Zs3MXE8jDO1Q52oi68u7PI2ttb8LaVYdvt+eCIoAs5EF5ATylnxiwuc5pvw8lU1a96
1Yp5I+Hd6v2an/7MGuwC81RsJFdXFTB6D9vNW1ReJS54Ohrao/2+MfoU/p12VAB994KNRopPUrCN
sn/2uLQog3nsAk5tAeiqePSs8RJxjid88jBZIrAmY7LvUgGxYOlhtGMJjhcWovCmHgRbc45CtrKD
iCMr3A1t622d5vge7iCoBEG3wPz9bX0Qw23EQ8M+efOXGNtewYOOZzowwZ60Q/0wV/erw/KO8Rak
LUAh8726FN9rq6PUoGZLzWGDqsjbrY/3XG5iylSkrrbwDjerHSCPszl/elwhb8CCBzjbH+q6a3c3
qiqP63CzIGpDIDKoJmznwFHOiuvFt4l+I7xdV79nqDqtx8zg5WQKRxx4cuWaeYx8LywCYHChgUQM
x0gmdW7N30HmPQKFy4HudVYoC/pOAIUl4BAchI0rs7J0JYJtiWJ07nH++acj5f0ZvnFFoZeRgTkt
4l0SBVbg79hB8o5gXYm9cxYAjMM6UZLikLgxTb1CFMoboon0DoNbSjfkjmuwfnoAQOAC6jWjOjoe
9FlUjZLDmXn09yXRHefjDTRCyMLghnOkTvqtPlKsv3ns8WjECq/kMcBqTUXHE9y9RzsctuevFII7
YSUdDB2vxQ3g+0VRobTk8I6qoWRKyYnFfreGy3rbqixkwoObHTEmylZtly0+iri5GIVRBMup4GK+
39BXLPO0xO8Pa2AmMH0u/eEkwKnFWac9qFLIr5eZoQrrW6rrRX8iGXPoPPcZnPP9ayG2EHtOkHWV
EOuLz4Nssm5b1E1WO+wMm2njmyKMC4et96oDbFS/8RkaqkOgmej99CqlJ1fvgim0591dgWNXgUIN
UBSGPgvJd5jpetLZdru2GdZNmEYGCbdYpQW3loGmTC6Qnsor/naTR7Nth+/ETohemjw+TaSQChqj
uaZ8MLDH+dUDbz207A5rHYLSgwblqHDBz/V24Cn17rOCq7Iz0DV6dOcoSp958uCUMrBsh32R1KxQ
nIIQLg6wjhVSBpJIlJ3Cid0IUk8rprcTuQAw0rNhouSxphFCXuRQwpAQvQFXbb6C2k2GrES1QCd6
uej6aX7CN50G9+PH6n/y9Fngek4vUvZiHH3GksZK4eA6txkQVmr+DGSMcouy51vfSPG2KF2O+xEG
MYLmgiq0LqmWaCpAnHyMw1wTEDhIa6+e5QvSyhxO0KgCDbkCq73kG9MUt0YVJ9mWzigJus/QPM/l
9zK/dtGEtP7VpII03tM8cGPFduZnUseISVbNHhTvJiW68f6EL3eOqkam7JLcnJSSCDMMv6cFh1dH
6lL3CctpsavTZeWxzmJhLGNxhDNSRarSyz29apU+DYOWpYI5ygJOTytSBUhwpYET1/94lbL9jD7y
QJtQCTDDrqWRMsCXKycvBVTf3W63HZo6RvmhBi98X6uxv83WQPg2wBAzBKwlBBLXtohLC/MrGzxn
Z5Dbr9Hs/Kwdia5jiX7cYL0g/66wJwHTqxkGUH+K8/SS9Rqo1HVf7ddzPAhvonZJA0YCcsvGMEQ7
BXZjETD1sAxeBeAeJcLKWWXqvdu5/le3FPL8Rd6a6T4e9zEkzNHdYMlJA8LBW65nYtM6h9aq9ie4
arVnSx00ypBvPPTdtoo9YaTv9Q16tcd6sMEQlAC37hQb15pCjs0r5KCnQgACRuQmjd/YFr/tojng
qBLxLa+hh/WBcY4FNtC/poaJTDY6/9PyxNwRiANKKUVuW3+AkILY7zKdqlHxPjDfiVHOn9P323IW
nnsCru2xpezZ8pGzURCav9a0VkpIDsgcWwL7bkUtkTEkw1ODbyWDlxg4T7p3b7HzwBtC/Ff4k5JO
1J7l14tMP2i6tFPlsOWogkB/5wKRqnOi6j7nHMqhLmUu8zgrH8y1y0X1u8w9vKumZlEJreYJr20Z
jKdO1EtnKWYIg34qjOm3phPJE8P9DVoNI6bm2bGJ7pbpjljomRFXz/u75hqh1gaPNvqqzfY9D0Lk
nsjS5m8WRaJhuCIyX/cjDKxS96AuxcAhQtHNyYxLwLZJamdQkWApZM9sdBeuyrmxiPy4lr7Jp+wI
1bsx2HWN4UWkdmXstBHv/rryPzQF0ZLRvGnK3Dp95EtDANs+u1KRdBCpxM9uFwnKL4dpHthuWbSt
vZ7NFA4BTettmAR+w1MER5i1+QM+oRWjji/lL9owpBPDKk50XsCl7xTPyQ73dt56aTmQEktUd0JK
AQmmPkVghQoInH4pBnlD1jKXP/1p6k5+Txjc8uP2B3QWVf+oGFY2Ww0uBuGeY/WZRSn5rRN+sUT8
2IfXPjrsIOp5pfpvWZ1XrXDMVKfcMvTgz9W0wn2UDwH4QZSRFDUolbqfWGvgN1n66ty9+MflicIw
LvL7m6orO64kW6DJp8pKgjSu/exRBNFg4TLFwJuWRw5kCR8tx72be86ducXhjGXvaNYleJzfhd3p
OjpSgvRy0d5WjsZwobfn6lY5Ub+WDxmeCeNVbMTUW7UARpuhln9fD0G7+Jc4ymC0axNz44ZVwoio
3McBgC2pdX4TM8IaHQf2LV0Xn2mzbMwfLC7SLM9c9UpIryFlBTb7XmHXVivoklyeIr2z16+niV2M
WDjKemyIwET8jXGyvt5+hU4riplPTkZUHZS1A/Ieo03YO5OiQQBe34RW515Y7DO8a/nTjcDiga8s
aIgq/7B12wJ2nEXFdzI9ltCa/xEGg1wN1AkUoJLv80NzkY2QH8xJ2NMgVnNLLCjb0YY7PZJb81AR
+LHQFhWEfimXwrkshKFravHuBDcG44mlLEjdjMPJqSBypBA0AilWaJtYuk6nr797E0zGip56mC09
FxMT4s90/4pAuRUzBAlLicL7aUe6w+LbqELb/wNwCVlrzIuogFHN424YGg2NSDABJttV5oWar6wm
mBwQF1ObzmctYsK79C3DmyGqpXLSZr3ehTKX5myMvi77UJ6ntWWYLYnl6do42IbgeV4/bLoh8M9d
LfnSedcBYSTlGg8sPfG5mYNNXl4gxTQ4y/nKmL8oisHjjWgqgtixVjb07oSreQdFKVpuXjyyzb+r
n8+nrlJ8Y1kRyawgLD1SvrMIcIXP36YaVI1lDfKDfe6iI/dd3cOb0H73uaCNlosyYsA6mzET+m3F
tLRUNV/xJSFZZQexW182N9OdapIIoCay2bx7VIg56frAUvlsZi6avyZNaPeZlAkna6ELNnMrP++y
JGJuaOKWqkZ3CNttln8JUt4LMeK9Mps3sbGTZJi0V4yOMV9fohbV6ikyyDn8963vq4DRENJLprC6
88aWIJ74AndJBkUEh7Q/N8ZcEvYDu5RJWDxFwUTh/P8dxYA3akoDstti+3x2Tq5i36Yt3q790JSy
WRKTto5Mknc1Wf4stFkF09qs/FNbZnglqfgVT3gD9VLOeAcHMceRLSdTETpfn0/jeHi4CXskr9Xy
XajO4j6Em4lKwnrB9NDaS1kAG+q7XcWAg5eM3knoC5r3CfrdTTXqg9iYF0ybn/Rb/F5Z+JdQtf+P
QEG/G3fYVYwNipGCPLGSd9dKfvrKSioAOwXskWb7yO/oL/1Mf/lMy1Pgykqt/qy6rjMcgegXBB3+
Q6lEooODOtfbiLQyG5mASYUo1G3t1KxQ6XE0Z8RhF0PvGp16qgT01ld6TLrluyIFRBedppYPSfEo
9lRJpgmZMn9ruXcV6XRqMS8YUrmSsK8twUbZ1eUW8ptdFaqNsEc8KTWTC9AR4njAKXizlkb9nnPp
jXgHs0Q1QxyjPyDxuCWZxDtDbm5DZipDXQDMkLz37RkmWUkd+UdOlR4o6sbLmOlvdyBrpwOXDo1q
O34Q72ZLreLHnW2AgVaTr8AFjL+qR8gyBJOVp+rVNGdIMNGrHDfd51fMbHnSdXU1BVqaFjgOsbL9
7C0aqepePSan0KacXb8KzS9QgcONvsgk4jYknQhsRuSSETIVcSmdAfaqOcXY+CqgdYYheKNFq6qz
91xASvY828+MIARCuzef4XqSWVoRFG4aQt7JsTYSi8tre86U7BGLvawimIEoLhvke3zRXbD4WH+V
sMvDbx1GkrwndFaja5sRYqd0lP3WOGpQqziKwRdAAZIqvhDCW4wXwln61usWmP/MwnObSF4T8Qen
TzC0rcBS0RTByj1ZgpCQenx4lb1uqnJAQWDF8Ekc3DquC6HxsSLqblC4xaZpJzF0YnB+3mE5SqiS
gVZ9ZaUIbZSxne2+yTpp/UwJ5rceiBEJ1hlM0lMyyK/75odm3t7LHXn8Sfvr8q9zSkoo65OY+fwh
vYtnm5VJmzxDn3VmlI96vYnwbdTVzZA5p5xs0d9RtUloB8dT+YCcaB0cs1r7WJ5vAHqoiU4qXzyT
n7Vsa+ebpVfn8bsTKE8bGDwoJ9TFEWRaLoWFg2P2X1zapQoqjBe0mwjaAjJrMeYiKvPmMWccxEOp
Y3OBc6PP7gUUWfAEAg2nPN32afmxfqEiADdMTC2WEcaPWX3WeL5bmApeXhYMwoTTMyP0EGQwSSCR
vzK1dXXeXVnBykWrf4XNIrL25j0ahG9vh9ERQTflEiwjFo+7Zy1wOyKgMrwns5N0C9hxPAhPF+hD
c6PmojKud5KEwoj585de9zI3CX36NUt6UPD0nwlvHTh6eHn9+8Q2fSZjp7gW3TaNYiVOTj25qiQG
ITogA9dwWEbzNIAcqm/LYlEekg9KeFppltezK0iFy8skwo+PDcGOHA0BkbIgedEtXgIH9q/H1Ynf
jyByWcn9vfl1Y0cPjo6IWsL7zj+GxRo6dlaTQZ26O+HR6s6T4ePCDTQZUd1yMQGWUrl5D3lRmhJ0
3zHXMNo4BNJnIbdejZtHWe5zn37yR2c3CObGWco9excJpmZ4CxN+61/zcpOm7hUAyGbSWPEglvDq
s4Tmuf2Cb3v1YmZgp8+fBJcL1S7qgdVmVIxKmGfdYhuXwH32oyjMxQLGTV6CzdUE1raWc77lOeEk
UNrvG9amiZe1kYKl3iBpgROE/C7PAMbvVn5Z1O5E4NJaSWIRLazDfL4Mk4J3gQEnylse4LvG48Gw
QgART0xg+AUzFnZs6+NjKpyQG6i8P4Dmj04yG+cxbqC+WqIyy+N+azC3869BSGcQaQL///XL2UV3
f3vd+FO5IuPUAtg0blVRxwi8wPPMZ5I9mIQdQQq56qksmG9CiB4fXYkvW4utCgP2ZS4m8QGYdBoO
hZcL1ErLb6oEhUbQrWQADOeSTvhPD0LT62gM8Do0BYGskPU7NVSeSSUnmFN9PLBhq6WDXoxqB8zw
WdwMO7Nbx8RnWNJWwVvo9sQsvQrRc11CeILmlMeUP3LUu8woSjpVLikR9od7uvX705dYTrmP62Ev
aDmFxz2U3KIahESsaPF2Q2DGB203mMNAc+vguEDq6TvE5oqhtiHh6VP4ka1/3LtRTLtpzTIQ0bLG
PMt7k/6+evm4SGfEKyBpKoIFKNzI70Hm/XkncfesK660tb6IRLECJcxARa8eYyA7WoCi2R2Rw3rL
Bjt9rTDpHo5WlX/sPx6EniKMhFsxYagK9KOBVlHHHy/EPySPQF+TInoDJb92dVKL4Cnf3qEcLFUy
OWztGmmT4CRavX1JX6NadH/mn4mMXHjMnDd68r4RJmpspVmDlZ8Ax+T+CwPjoMRFXGBQgtcaFjgg
0ShLompfdUZE4diKZlKnIKoCZ7WYeWSig4tKmxe4sJEkIa8tj1E2LGmq5w65Ri92bE3Xuk51Q+Db
xJ8EsOAkll08L0pLplxKMj6DOnG9jC6AfCV9pTv1YvrrH0wIs+TzDRWSVfn6jdk1TqN9ezLUd8y1
5YrQ80Q94gpvTqZCOfIazSLGvdXD/oTXkGbGuI8tEeKCkNf0U6jrp6cWLjZHoYBw3wKi3g2AIr3v
kNXYGTQu9DMWT887vbxUfVF6M3J7bC6/23dxXLyIEM6JQtzvG/ClLzY5+RMts1pu6isJpkTZHbmd
NSVGCrE9f7kZZ2TheGmmKnKs6GmqlEK/w+HIHQ3hhquoGQFsqsG6/fmWN1I+Uqlir0OrvTl9v28h
8priR9ZgXog3h4fLItdJwoTWLU55zI8kFPl5fxobEPc43DzIm5NPk07FaSkbXE9rUIcfj7KFDRtD
DxhzVi2daC/zLxXYAokxsGMrwnmfheFG/hHN9Yb+/LoDVAgBUqYXiJhIHYqf1cn0V+cLDQkrqLhP
h2rWDIvFNx2/OhdjOWODY4cUg4mtR6b0tFF/ldv6M/u8QYjvv6Fgnm/8gmGMK72lFkCnKe4Qs/Dk
rLqM1gm7jaGKbS0Q4eJ0aH3KU6XZPJ00FJpXpvz/o7lZ3uts9ADqOdmDykrZDg17h+eWHPXOapFb
cuLBE9+uOLmdCnW02yDP9rJkDFLnmrrwbD4bjFCF9MEtu9Zo/s2X+AX+CdEreG34CAUV9EIUCJeL
vH8Sx5hgnjxiZ9qwqTqsBOA503t/6eRh2UQP9ItAmTsVRHxkuvlVa6BYIC264Vmthr/fFZzZCqG7
uScv8cCRHSrVFP0vq3PY5yAriofP1Sx/cIyH8SstaLVnQ35xwWsnIID+zyVhEaYD0ba6t+MPo+td
1lomGo06ko4mpzqnKgCMx7PcTZyH3ouHjMvavd1rO2alrwwgvOfVHLtQdlQudA3rz2FlOowkeMcY
nwXnbF5Ah7UbMT2OT4ESMPd15RpiHVRHnXsiw/s2id4psyZn3/FfOgDHHpBDBDh2u9U44H6oXvIH
4R60zvZBcEQaiChUvRXPjKpscg4gjjE8E3nRutm/pUUZTdfavbmt+wKfwV//l838vSCXs5+3o+R8
Y0zD5cNsX8P6wYIooP9Qdu+/AFYA2fVTu1dokM11ckA1GK+0QznjV23dxNUT0reNqvgVpoVU3H5H
R6TfKdOrbKEwHl+q1CXhUU4t2HRKola0cHUvHonmOBOA+BQyxy8AarHR7d63OdZaEKqvgVaMcGYQ
xdYvcfTEzT3cfQ4ofBmG7mtlhdZFrv0QWpHhs5oe9QI5nAtwx/k3jYei00Sf7+KkuZ6VsVEAXxAO
HU2OHKBLkXueQZShQ4+VjZV5H8t7xs7bW8aFxiuGBpPhwBTXWhEEzW9GSkMtnm6xSXwfT5ObzrCQ
9zQHgYJsOICR1jom+FLFhZ5K1wJsnz7nPggIJjUGaQUyrI6HNRJ90VDEkJGuaQsRCTv/LijTwYN/
P0WIlGREw/DUDltqFWgFaKY1xFOehEMCU3b/5AP7ldjb9tBmlD+RPzXy2/xhVeRDBhlK+n6iD/Nn
rWkpxCIllNo8IAXKQcUiRsDZzhYTyO/bMPkMnD2PUFL77R58eSnt4zwKd0LU83DL+lWBJgl4E9ss
CkhdC3csUofv6msE7VElvWMgJYZTcE+Nd9Or+1tGNcBLLcsOvK7lnknkwX9r+zbf16Rlx4Z5tjPT
jw+C6MapWZdeD71OrxA9klPr1FrwmH6s1nf6cvI90DW0j+uwzXHjVDl3A2iqj6j6jX2tUgdFcCAJ
8B3nuIYUba/yV6cnAVRKu52j77o/3cxpvQQBn/uhZ4sywWZqhiYcP9tREGL/zcSHzI0cc+wS2u8N
tL6v3YDdSfBDciXqdyB2JdcUwEOhGm5FIsEdHxHwh9yYZ5/WQlp1SEZ6XS9ZIKpAQxlapwx7flKw
RVA9DiyO5yGwpWanDTA3pXdnSVtaXjxXYsjFHxy1zWHsjMFFbpbmhNJlEaIorxn9vENYL5+Iq9dn
H1coR+UZkVcDiR8ANxI3TyZOgKj2MyYXjMN1ZynzfulUrW4c3fGj99NQReklakxUUycDQq8+JcoM
GFgDTCU6Y1LNL6gKAY0g5nedZoptNJnExUBTe/2y0QQM4qCSW5Yd6WGyyG1GOl5Ib/t3834LJ/mV
VYgJSTsQBeQ5FphioGv+TOXIG6ISKr+rVOPmsYmjjhPU4zNi6ZzdEqXHT79hxwrBkRKw9VZdGSM9
w5+o+cM8zJiFhc5EPQ0KbSLRdnuwTQFYOnosZlK7a6uxXa8afd7UuqTVS4NllPHvfEnYONiO35fO
C+SFs58gunkXErNVFxwaVYm+dtPkvY01vuj+Y5MN38Q9flwbx1l+VbKmFBiKcepUJ8B4LpmujkFC
Q5uOUva3AYduxRYCxwNCz7BeY6oz96sn7Q/BAUKQX/nXw08g8zlng15B5ItxWGdcqGa2fYnEbyIC
v+Hh8rScGvsR+vNpyAVmzEnlYPuuD0fjCXsZ8ksQGLXKVWQYqorExOonJXD5MrI1INBxpYbYyJix
AGY/vdLizZlXca8D7BlTH4w1Cj0/Ez3DijeUfURDb+1iowPaeB6/9mBB9SXqu21BQxd7fNZaTPn3
pMTci+8Gr0lITYleh+IlK6uFUQzStx2yKlTu88yS4V//IEP3xhKzqYAsrMvMRD3WWlSVHJqGNfMH
BLnzz/j+Ll8suDEBclr9ZhWRz+htA9ALlwwjRIZWrpVAmjECCbiKeyW665XNj43su3pZw1SBOeeV
TaX8JaVTTfDMTETMqsXZNy/cDCw6yLvisHzrRS1oYLhca5vuMFu17kcjL+qhhF1ttNRYRQp1TsgO
GPlUaQ1yFGsANUTJy6YggdcKN6yzra8SQu8tv2L7X1arjDjcqtQjsWMIUMmMF+X9vNDVen3uGZb1
Ubb2FcVdguqEl847lUYZ0ar+GykzYKRARITFkcJCXXPWr5iIMURCrdDx/u1LySVk2LxeSOvWCrJI
QIccQ5eiL9lltzvbjIhU65vVHZ/CI4kacNHCiBN5cY43CLBYekQeAV/C3d85NhA4AE5kHblhzFH+
cVrBbBhtppTfpQ/6PE7lDOfYlNcXgR05VgwmZFAARe6hkmkcvXSMH7N40Nm9YRYmvjxFdAujqfAz
rBvOkDs51nulJiP2/QSyhbfHlzHvmhm8Q+HEt8GW/b4JXlMLFJUy5lM6hU/7pTapHclPaFq9nEF5
JDb8/I5DbgwTtaSWj6EcKJq9tu64gHJQLLqvIV4GzP30a2g9i881C5mhRW5siMQsvozxtjYZNHa8
hGIoZLiXpqr4QcwLaI5p8i7fLUq+c3B//vYefskf2pu1ovQWnmpIKCtFa2JpzCYhJBzmNs5uY/B4
uHaJnyxTfzKHATpqg361D5WpFt7tdIkkeLOKYJAe5uFOhB8iNndAMXj2u5WO9jDpEjQaHcSZhsnV
OlHzC3n2JZAeC2XkMUH0H51ygxgKtjek2yIpWSvhzNu/GL+4qvyROL+q4ZFHu86F0e8/tqEn0EXO
nZoHpBjPS0bnQYV8cpqa3p/WYyE0aaytTRXyWFJlbWxH6rCOMl03/Jg6eTJGfOZgFL60POG9gLyG
CQCytDNMCkW4KWdYFtyvWOTuZlPnVhdMAv0HA7MBL0zeGKHDQfUB8LEfrZVkg4jZVYeBDtmvI0NK
NY2Lc4SvJk0VKQVnrhdUgpnqbHV50RizCG2wmN3ybdQ1k6LWPDY8AoWFxmD4H10SGy0fM2UGLmgI
0gsMgYYIER0myJ9AAM1yxx+sUuiPsCRiNO+LofnChFTX6eF6DHz7RlY+rd4PTSURYzrCVCBtZ6Zi
eshgcnMh2CjlNXVCwv8jVWiGaP6oUmBQxm76UiuFVcH4eDYnjWijY5Tw6l6tcaFiFPyb+fXVx0PG
YhduzipBA3RChJ7bFmKReKmKzYfk3LhZTiUCmrSZLn4qmqmuchYOzS+l44s06EXy+UIsCqqhTJAT
SvAZ6zebkMVKHH0lU8n5iEXqPUKgnS8V39fWYhW2I2/ZYxhwRfOIPnRse5rNo10Qq8RlbniOEraM
X0xjWOaIxRpcnHvO9cqV9pioxtntK3IRS2Y9WCGAYR9nnORQD5HUM1RH3G8lsDvAbON53nDcJvHX
HmQr4reOpthmsYnhMllDbXc+VM0txZzMdEm2W0PnVEiQOrQ47iG9ZK8J2qhuRPOdXKT7flnto5kR
oJu4yfWu1B8qclIa74YYO8rep2Av7aQ5nM931haiPGzvvR1VrVLz82upVk6YCISb5iTQvqwcWJEb
fOK/tsF1BMr1gRoNbwbp8TtLNZm6C0DI9KgEsYyMPWEhU1RuPN37tm3MTOpdwCdQ8YcS7P32Jag8
I8qU/eM9jd5bsWOgSvTJ4Ig5MBlVxtg6WoDMpL3hk+jYOB/LEKFzsthce5FHZEpqEvHhAJpa4+/u
Rn0RZbi4JMBuZ6c9xDW87jogF93ZRTKY7I6BsHquqaC9WpBeZ7N1eLDW4PG8zFkM7cyIzjcE4XTS
QUleBCSMkKKANMhm7Os7ZpZY1r0rPjnaTeivAkTdUOrkDLgbZDAlVViKHUOBiE1zMMHSKPCAY861
S6TrWaGdphHnrlq34evUN0/Wp214P+sWGNogEwQq/5mHFXriLRFkIZ3nOkcQZWbYUcjIb0ywLR2J
KAMEbBCRi1Zeh1BuLYmcLC8qtqjE6SiScmVjj7Enb57AorKWPWwOWSgXgl42WjHzsNchxERXN3eQ
xWWXCfcNg+9M1ryb9WQX1o62YxhKWGCykU6ofMf4EhJTHGDFh/bpPImlBjgHv0lHlDhokbS4dPrG
fTLy2M2Il/IU/zXnxbNJcSQ7Xk94bI5y1WXAc71Wrmu36qt880m4F07EOvBUoBFfVVSxoE9WXvpP
o59oPuyKK7cAzh15NFjzvHp0wts9O6zCITcVaPMVSnWymUy59XrQVGUX4QbslyZxqm4fhC6JA0QR
Nu5kgvVipUlUyGSdJYMJ5ktg1g+btVjuB7qRJfjHDxZMN0bOn1a/QSG6UHOugGckHpNNSUo9oi3J
McthKJeiF0Nmlk/COcZu/RlpBnYEjDK6w5zSM0J7wozemlK+zUr3G5tz9t/mKqfEFR8aawPfo4XC
mAPOvzrl0W/eyNZ338NwZo753w4qGjAoaPVlZJSovhPWvVZ+Z31LTLL+YKjiqo1jEdm824JWoXVa
7V3+tKMQPaXcHgBCHHh4uFA2Gd91+Vbwg8OgKV2jRQ/rGfdpSs81TLc7/ieCjFe/+aQs2VT1ddMB
VuxwqERbwEiY7BJwh1RaU5M31masJIKCz0lgIV8+7WDOvnwChypfkSdUjPLkAM0WbkFA1mK0Er76
YgAaGMccpMk0czSDL8TBK0QwnBRv5U78h8xU7eKzUB4VtvmY1HPiJ3S4NQvzbSp+4Syy8K/42V5f
sbP00d49tBCy/YcDPK79gtVSaIDYqA0G9Fokdx0DqP5zkJ3wOiLsuHexckdRMFAVOmzkgnI5sWf2
qZHDHbkQsdK+xmDc09jyui+068iImsuPfgnpHwEta458bJphsz7lkniVzbYY564KDIqkTE0Cvy75
94/blKEcHN53/2m2WtUV6/XwKTNiMQ2E/Nlbwtf/zxkhIoKY2oXU8q1aCrGconzK1N6pGcUE2XcL
JTG+P75ggZldOAYPtG6MOjzByFgPRNaRGNzS0mwQJVuapd10ZSHfQJeqgdA/8wUvPzXTFqeqOqu2
HqYK+u5w+XNqp0aDFmmGgcHhVn76Qx414s/V6TVPvJrqqwp0YEFloe6NXmmQuP0i/+PrkRFPVPyo
X9tN17oOLaFEHuoXMLHAkCoL1vO5pBrh7cJ26+Hc1u56Fl70wGs09ovE8l6WWjA3a5qOMtbOw9vQ
rjwDl6hUGZNWz46F3K4m0BQmTmjcA6lK15b6aj7oKtR6gtfvVgnOj+KCTrLTUjHX0noCAp7WpT+s
reKz6SCZW4gANjbjjEt2gsNoOgzHpb6l79ekds6VbacSa5vxfaZVtZ1q2Q5zCL6czW7wh79eVxuc
p9NzjGm+9tNpvyJWP/IltH35Z9V0ouiwic2a4mZPHMorx1CBLuRxulTh/v2ZWdHcLzM49zx6h/2L
TwPxW63tRSOKgMS9C/ypRFCMgi1DW7Y/LrXTnY1mmxZNDTZDZcayomGWM8oYhcdWIxQteABQLKb+
TJ6YbRdM4D5Aqax4dd9xcIPUNTm5OZ4oa7FGk7MnCtFBId/sUA3xzKeXbIph3bYvgq+EmtGRUKr3
IvKoYcIx6RAzIYEBtj4v/GxZIX8AxZsgyAZxyWTXmyOVwUCTLzG1b+bXT6Q3ZJBEuOdOsybVa9aG
sFD1/qjTkxgoxO9NnlJdvV1oYJsa2YX3dFZwx8JPsFRTMU4v+r4DIz2dMCBpgV8NQM2LXwUEyzm2
pUpbhzN0Zy3BzmHF3In4LaOhebhv3zM2guPbLhCv6oBS2QyID7ecTJVwf0cnAXrYu0hKknlBlkWI
c0VP9CANPf6EIfpqr8bye5c4IflLeRLpys5CL21Bo+qjDswjgoqcxZarHvEtE/ptWzvzggM1przu
Bo16bkilwuGNuNtwUgNHePvyZsFGBKRYAtZ9HsKdtH9UaGTuHYCald9ZHn+DDr24zEjpWWAMHwT9
hruAZS8DUagL6f01j7Ru1Bjm8Oyp4VmYf+KXYyezzF9AWjbsa7YLzLKC90ILRO/1cB1Qi9yPePMM
Pmk+H442tQGPeMwyZhltjBfjd8pWlp7RxjRy3GQYw9B1v/IheJdVq3nn8Pry4B0Ec/JZbAkeab8D
Bch5hoqOagy0zoV43dXh8iFFrXGXmpRMZvjXjZ3SuWVSD61iKbbCRaBIQK0Q9W6D50qPZWXviz7I
LpI3Yd9ND8bCXwF1wwVebrPb0JfxjjHGLhdur1qZKaj33s8TJk7MCTEZKtHHdgNoUDPYAIc6+cme
2YMUhItOx3DT+9WDor2gtxsDGCdnLrptRAs+mJeWTjlxL86SjgJHJwcfpzSyB2a1xvdLCBz3tWzk
QpP2xAdqYURmm9hWextg+scO85NdsnpYRmOQTLtxv8DjyCbv5otaKCQq0iir6yL/Bss7SDU5JPtG
HcHQc/ZtArEDgkd7tIMBt2Ey2QgPHfTWJxsv9L+56JrhR6MkJzLWZtCQUXS1s4O6kz5k8towsFUH
doIRzpTqJcPLqLFLPQetYCojHIBycbCsVDeWtJk37aMH7ZWxdMmr5LM9AGIEO1fL6NMrqgVab9iQ
RdVq6PZkDpwx6lJk2o30tU51HbJccnpZWpF9c9lLr3mgs/R9b9XD9rjGHcbqZoJliBlAdRAeLQn0
UlOn3KVUfLzrpQ5YXdo3ZHKzJRv0nh1oC6kX9wckDvvIEpMfpTaL2me0NQYpj/3FDcGwdnKYiKTU
0D9MOB4BML0aLlyV0gV9mljF4s4S+qMpPouYu6NX4qDXLvrduq/0WF68+b5XXKc+prS7XgU3pBEd
5HbsbxFyuc2LHc4J4B6mJzJ087hMozE0zZDo+mv0PFvSVBOxLAJb1+d5woQ7MJavBaYK9gHPVQ5Z
S2DUan8uXPPe7y/ezCKw/Qw3ml0CySJRVefBNsp0lwt2oDhD7TyIe0HghHJUk06wdXC+tDtyMy5L
rpuPE4+Q/eC4wtabT9S0DfwyyB3OlBpbzHdvYImoegzEIddCvlXF3wQD4q+T9b/wgovmKwZqbml3
7nJSbCEU/dbCVXKjwf08eQfiIYClN8HWtcXJafeEXw+S/X4Y8hvzKcpWtrki26i5sXb/jNn3hgre
oP9nFEP8wj9d9w60fQg4bqvU6tB29k5XVlXR7Ir/aQqyF9Es9lgjM2dxrBUH93iGqVngJEInf39m
jz0s56/B1tHlU3/q1IkaQonbyRfHyn+Rac/MMCC+ZexhK1tIlcvVcSTHyE/RwSCZMqI8GdMHw/0r
2QJmCrtQUz5/I/iUd65pJ3KOPxBP3skfynhlubQsISw1AQ+zD1XwieVxQni4wUsx9/oQmb+FEGfW
NWnt3EWgLD6Rzz+ijcgedi1Hw+CrElt/h14byTpTOQR5RQOx+dJ40Y6t+rca8Rd/jJHgvtis7cSt
nE/s/hSE3rMehkI4rqZV8JT5iqtVK0mTnN0aTQKvA30LIk8ucKlnyFM4E3hXJJQyD+MkG9QBHSl2
auwpnBwQq7oorABqt1XYcbG8Ugq/LB/7mgek+j7sFd5qQxGenlfeyl78I1vyVWs14YP/ktpJyCvL
980cTxjQ1I7XfWAxA5muhWAgfJyaK0u66etuRFOGURe1TNyTJXxDuVhdKnXnYNOsybQjz5a95X8N
H4pVS2F9NMealzDX5ZLYsPbCscF/A5WiROpJxJc450hIdLXWEZIa5Z4AU8ZDcxl/03NSX/29pLk5
5uG2Ku37CbLmaQ4Za53PqNyf8yYAhSW3a/uxeT/5GFXcMjSrji2mMTBU2QpQAUrwf9gMQMZ21Lfk
N2mHsjzBxX3SWMHmMeOvn8ZwNfNzExbatZytrLMhpJsuZP95wdPpQVCJ7GP1iN9XUt9eRcrKxl5n
1YFDg/7skMd+IX3oHZFAAW1gH6sVi7ANP40jySKIOstj2LxKEa4Iq4iF8CjpyeloYJsKSrS9511m
lHLP22mN/TTyLrWk92v6If9ZaHSh/lL3p0xWtl9K21gruJ5S6us7VppZAoitg1MbOzLeHQibA0nV
DjbAYXm3y/cM1HmzemFupREjNlDsC0j2J+z+Rlun6uhonbNBN03EcE2mGl5RmXPA/WBYsIFUjGFD
D15rPE2AXcghG4GUQrO/VmNjhhPMC7I85NfDU6gDevw4jJ/tmZcdBR8jIzlSPGsPP1K2gi8yz21P
uovPQEH1ffxs9RnfxUtibHp3KcLa4gWXgBowp2QnZhjmm3fd/VVW1SKQXSZOl8RLfXwYskIOCS41
a3Y0arzbB2g+IRdEvwQbK64pNI2YP81MsAJM7anlbrNQ8PdQgLv9Z5z7P7RouoN5N5AEMjG5VJLu
logxkGFXe3ZH3gddSM76Zb1T6030QE3SiIMWic6i5KM40awQkR+zprvWBWN5YDLKc+PE6AfWJuqK
Pio/XziJJ/GeR7eGo4T4+YtPeqg7+oAPvDXg15HhCm50SsZbwFZHYC9TTTi1YQIsNRTBEIG8+LX/
yBO/j/589+mU50E9lNYw+YUTmp6m4Qvccav7tK1rxDkLZ6kHmVGP0+Rm/AndWN6hKudgIY2V5I0N
R1YaNCQKCdLB12c0wZNZsh9PmRN4xzQpsUsZJqAObbNjBLiII0bFpLCsn+BvawWNuXEW3j2BCjx6
nAZbSEQDacLkGVqcaXz5Y13Nq1u9zwgKw3YeXpTu2NTMJhwUKlWN9xR68lK42Q6Ki9Zu1r0jV9yU
YL0O1+MkT72Of5cVKeeeBzhZQYZQloQbmAQ/vBkyULr00XYZdMHMznHozAH5DWMTZrd0lhY3oIeV
Yw3DFAxPd3cDMDMI4d/19CE3o2wM+eNOw1JesqByEBA7O2bpqFPHRP24inl0r19dxYNXPivh5DGI
DOCYghgl0TpsJIWCGX5mjlWK97lOMxYQs64Ehno+7qBE3asWRvT5gR3fUBhWne+7z6Tqtx6SZna/
YgDz4w8oyywe1uHXa5K9Zhqqqyri1TDE/sa+Q3EsmwtfO5kuzdogqK+pVshhoZQyDLWhTpbTYrhO
Z9wRiu/Zq2QHeZrekxjo7+UWMC3TlkphZR8YxEvV67xM8Yx/fhvCicQ52Tcj9tCGsV2Dp57QNiao
eutoFkFxTQDpFVPVs83zXPUZlA2SMffMxgKfDKVMZ4R3n+H13fGZihTC/A7FYookgcH5rbdxKZok
2o4b/pH+ZKbweFzzpZjGlHe5BuaUDGJD2/ZM54Ibya0Sw8Lu3z0KIGmh333J+g9vLvFUg7dR1OmS
PNLeqM7bnYFvOb/H6EVLbp3d5cTdZmFrI0UGk41UhqnfSPA2z0wvVg4KV9Nlu2/4UBsM6HvFIT+T
l1t/XD85VO7IoPrwl6CjBPUxMImeDisWArbdxrIPT1MdVK6qjQtGj5FclJt2NlBEoJQLHRuGcy6F
QK7LYgXHeeAsRsGspLrebYDL2+icinzVQVtvUSbD00+D8JpJQBGX+PcgF3ctU7AbjHaPk1xcDSnD
J52ZSlgBeYeQPeu9oPn978HwX0uv+KvjFZ8nn5aib9ZjnSHa0VrYvjzlDuC8unq78h+4MgG+MDym
Wa35m29pJac20CEdCgQiEGmog8CDwxWxnPEp7eFwQ9uCiXiFn3UAg3yzSb5zrwe8EOGwbUnkrPlM
kwFFV7mXaJezlDrjqHhZYi2QJu8clHo8fTdgSISOp8iJNiuwFdDM2JWgmInPVIiDLTbJVC1UDgjl
/EV8wwbz3begYfz03+2h1amRzXEZRMWqMAUdIQDOi+x7DxDyNEm8zIGgNwJL+QqjyRwlEMGbl8tE
ivP7liqC/1/CaKygsHDxi7DwsNxfWz9S317RyoaE0zt+pX7CqHWsVkdUGQPMmetlIVDPA69b/BZa
mbFLtHOj/M3v7Y235YzK9AhujBvvQxeLun3WiBBC6xXkMB3bl61MX2oLQ2EjQf4kYBCvCFOFnll8
5Ll6BQubH2OI10/woOq7Us0xqv4rk6UBfJZJ9p+00pBrZ9xf/hrTZNbm0bSl/dPhJI3bEJDrvg3b
pGeN9MPcAIyg6D1pgYzuUi7E9fsBCLu5XBpqPPX9D2crbZw8E8deEgcTFeyQhqIgBj8KZmTgzoJe
asYA/5DKYjR0zJ6XkZZpDf4GJ1M6xDfTOwjYJgJksFNtbwRWpXu76IJm7qnSgqNn9OMi6+LDBMGw
QzEu5DGSx6Ps7ubiZueDsO4kMny0aR1L2gZdGnwdupC75bCFJgfGFDn+9L8EnWx2ixCZSCAprail
/PPQmKYc3zz+cLzxY6bkGKdUAc5bQGN7F9+3wry3T2BipONLkGanbKalgFAOgMc11g/BNVxjGb41
eRv/JpvAm3p3ZdesE/1S4XbWlrSIs/i8zwUkWdj1x2+kCK+SSIZA7UCl8E0ojp6G0XjWHATAeSLo
T8vOmf2KPEouPyk7VlWRefioMQ1myh9fHiAWJZ92YLSKaa9x3faTeY6DUGNhJ+06B+nB3lnzNg7z
zDgM9lOmoBBp7svPF/jWktzeFxeR4BRYxBwL+opV+W0896Vb6SMNEF4LSHBad00rRCta5WAjQ0Lb
LuGDf+vhqryLrq4I6c1ZspWcQ8U3PsIRSwIJ2nwUXJdKdhGY/VQo+kQKZRIhJLmOInZyEZdynHgL
4SlaWPW1irdj65uCwLcMxuQ8Hvef55m5Nrwo24aQ2OMy05/keOQW+xUywfynMEsO2XoLfvzryoZm
u3Gmv7qlYdfE0hRIUhpkwT22DzCmdWTDJLp8ULtbBo6Q2Ryen+iUGR90tbtj/22kELloT6pLpmF+
eCNRh24M4Kf98XMPuWc6Gx6MbdQ1YyA8IsjD0Md9L6K7oC/ri96w8EYpyyoZ7DtgYlWUaY2X0G99
gUYiQRmZMYx3PMmiLfHGI5kKTlB/6UPLtb6kdUFneJDm7A/1OXmzAffDLe7/rMei8BCXkxma8uom
5Qi1u0a1BGjwybAomNt3Eh4SZk5mvExAXv/8w9HpJFfxPe3GUqIFWb0gLjfHVPYsuDgoLIdRQMZH
GzrHj2mLbgBIlQDJXttMVHN3IJ1dYwvvS+/WHlVl7DddKMFXiKCHz2yYz7f1sp5tpCPPW2xcMLcx
HkbEuxC3665m73835DQPzlAf844AA2RDwwJRV8Af2O2bv1HFjEbNeulZJCv+QCxGAYwhhkisM/pJ
XND7rdr7nvCLOV4qDnyjicc3j1SK5AKZaPgPYpj5ny6oThVyp4aeRsXg6dcuQ7ScYzx/kPxJYvbR
LDnuk7bYZkeqi5mRalqANhbueT3x+5D3CpJAk6XEUweg6AKqgKbVBZSw+wpdBGjr4FrbfiGcNQis
GQKgrTF/OZmJcyUB90PGXY06fGjhY/L2dvz277PxcYwixOKq0RCp4AcwM+zdH6lnSvFzgPOqj1E7
9cHHmITKSH9leWsFRpW/1ksN2gk8Sn4Itn7GFtHkTHkxShzkuJF351PrEovVV6uj8mQnAgOtybf2
gDQN+/gJSsYZmx5q2fEQoh3wWvAeVqdpYGhWCIy/g8hWQg6AekW2s1r3EpZVmsiKkL+BZgvchMnO
HUFlB8fmDIcrlLU8vvRyBs9RIdBFlz7YjfOp9OdOUOkD3ikqCknTgHmZUwxJ6Nur4xMsRiELXCM1
0rRB+vjRa3F9uWwgm6zhrSnGf9Ow0tIGgiYJfYDwYKBP/4IRzsIu27lyYwHZDwHHkxa+MJ9vSQ76
lEgUR8ajlgNLUiVbZ1mLNc6wpSFfVk5vHkoGZCG/LTw0djO6WfWWBcDV0l/GFC4ulAS6e1HEI1RH
ZS2eE15FE5YN2VPYZmC/TWqhStflq+8AIJ7NKKpV3wlg3efvZajPEKSc9lbNfxy3ZUo1TIcZl1x5
8RU4rNw/unC9B10T6awsV8DWue2+l0rFkq24snMpbCRHllj87UWckVVI6J7B+ym+SEoTA1ek39cp
CoMiahRSVzFnxZGGic7mubqRKdvnhJsGfTfWHsC/DgbiPRpsHJcoly41LDZOYZ3Vdw2MdSLMxSZn
Fnxx4nzsvl5jv6/eYwB0QRH8IbHs+GpLnaGOYOOOsM/Z2npRpcYrrWyO64NokdySuRbWhBUhpENL
43R/E+011MoEUZfMaKAyG8Rmzii6iiOCT9TeLxg5qX7/ofiPkuHXBzMFApd57fX5XHOPrbT8skNK
ITYEOMwyi/oOGOTu7KxUq+0LDHwEDySif7H6nM6HDDBNoLb00i+iSFbgN6pkxAg1QsrB+CfUlhfc
7/mcS/v5buEpWwpt4RsnMlMRL7ySx0C/njnsrZnR6dR+ZVyyW090gFBZ/nAxD+JZZBWYUl5wHpUu
bjtHMHK6YvTNARVCHL6hcH6pT9hGIYe7FRRlYHR6DaC/PlLJHx8ltY1HsJDwlvIJzaknuKodg5wB
34Lx01f4dN2tnRtRGcqOhF1EGUiLsRwKpCOHo0F3XmtzfezK0FlpDYXlserulJ/AiRs8etULmfHX
jTkHn8y5TncGolExBseJDCwjuKNc7/3b3LXNCiwOIzNt8UC8sR+U7UWKA9G8CE94XPD85EkvS2y/
B0CcwEf25pSKjY/1IW6dDB89llv4CSEoK3s8poizT3wunIXsEjDe3OTrXqCSQkmhbiHoeHm4duqX
/CUhM2wBe6AC65Y2av5YYPbtbnY4If10YUva+S6vj+1pfEcJjoIpymB3oQkhiWXUtvWaT2P8NNV3
49McWpwxKFFd430Yu//pcWdfyT9Xq1T+Yq4iTK+HQiH2CvHveGV3KRCoNnHqQDA2R/j0kL3ZN/ve
TRLteZ0xkdMdQ6LlvnJb0T4yDp+TK/brqwuDCpoWsZAnftyVF7iZB8A4aQ+GlqsjRzliSk7zBUYw
ycyBqnBEXxCK6XMM7p1BPm6B0HnAjbzCJyYUzhzBqPyy+0p2XpUtlfUbacDrEinOiG6MQZQI8KNF
8hLCLbBtA+zPplQt43NedZ36CwE58BR0WzWeQntHTIdDpNSaK9VLlMsSC/4gMB6rOkM2l6ZmB1V5
8K7zW7JkeV/Cca41POWeBlw4UU5/mCxBYVeVpEb8LEvFfdkbWpfkcYghxtrKQcXOKHVEBNRXpzhD
V5QZ5A7vJ2MyCrDvycopnlKQ0X+qyZoTaujKf+DRZnsXFMNwDf12CRolqbd7aQL7J226/RyzARya
eJ2K2S+qQ5QK9qNqvxp3H4Y+qw9iCPAQeWpp0ZDOk+jBb349/D7ItSAChyWFKbwJnPvdCjzPuyvC
NWmUqpYn0Tl4SjUlHtsg4y+TgFDcR2YEljO04aVGJKDVI9RrEJ9iiMRT0IH3lzRNCJD6tVMNjq9A
HYhIlOZ6bNpYkh9gccgTIc/ECSCP9K6PD/OXBAM04pYMBz4FyielQWJZNcGJH3eXMgq+SWZMpxBs
V8F99OmLCQONxMwTM2GNt1SfL0ddh7ZDyJy5I//Mj1NkxhsU/Kc5IurHqW1SmAYIcpto1UqFOuUZ
InWIHblijgfM52SYPOMb/YXns8uJxADn2xWsSCk4086lwTPyAwYPfGexn7yJLUVfTP7g4zNSjukp
s7+I2vjA5RXbW6/b6xc6CI44UhjR7OetYllOKraHFQL5uWQpbQK1dTlxFZTebd5od5icKf72wmOZ
Vb0fP70HjLsAiloH+vv8/VNU3hxc6brdf+2fvZstbz0ckp2ayU0dlURJ08IS/piQqPrByQ0/yrap
0XVcUdEjL/nz2NMC437ywNZ7YIAXSL+KMYJxsPbBef87+Yt8UdxglxT7ltkmiSO6FE/tqahhe5+F
M1hWCdWyazDAIff7/QGzz8YgP0wsLvQN0uBeDXkN8BJI4SfiyQnc52QmvxFHmxrnw+MfAgT5JuNR
Kg/yU2v2Z13uA/uqzLqCym6Vn7F3HrbxIXV0fexriOcRVutRm2CfhghfkvJqIBjwf/KT3D9Lh0UF
HmUoU5bQAGt8EcD+a7HD5h26TKztGAdLCYghxqEQS183eplRLOQDQ4zlR1J5tajIGwqq0wumazsS
ME4MAfA8+xnbOHUlW5pFVsWnm8pKJQ6pWOp4F2OvX09A3fwCLhkposRQhx37aHKo+sSDslEHZuAc
uPtDcxxfwotGPVaACpL1zpG6mpw4CD2cj7YbDoFPcyJ7boxDSu2exxz6K1CodQr/pwHH0g1yIRoZ
d8bH6fO8ZUo5y+WwrMidhCLfOCEEbIy+kI9d4cAfWY8W0uraC2j0/bR+qwxqn2qX1S4H1r6vD/aI
lHU83kxghl1yElMd0cJKbFbaz6Q0yH+6kwjV3EiRaRtY8VrxWh02nQR1rWsmGX0RjAr3OmlcgPbo
CdcXeSuvGLLFGRu6Mq6kKXYuak3/RicM2azCNE3GZGI4KGqigVkRJO7ezpo/RuSZp7fKLGU9kBRu
il9Omi/Oy8WqsH94cbjuicSWwr6EzGouoM2S3RfP9J9x+p8AwmtKMl5z+ims+iq92opKMKhI2KU0
nK6K1wKIAWu0zhHZbqOPA5EnwlUAQMxFzSMDhPqe5g5N4D3Rz3VRl9cy1uuAennF8NCAJ+IKosc/
txrqWMxBOE1sNOBDwhvc4BoknhSIUlfir/5mQIy2g1X0AQH25NLw2wWPMGw3A1et7mYQtsaSWVfd
Vp21Q00T4w9R7ZU22QE88njeP50u754XIlXGDgEVQHuPTfR7H1F84iG1MckrUxmia4ewxLFvWEPa
AQBJUCJTfC+5CvTe1yaCbg3Q3XfKv6xoJawnUCXvcFd11Xha5VeIQXoLVK325HjJIf3chsejDxQ+
MhcvzFpy83KCI1xT+YfQYT5hLXKC9ivMmRnESnPVTCrWysl0cMk54Txt8POj+cTZooBJHIx+tR7S
ZviSBVfLvUIVuNhnZWLtdHbY/th8RAvrQr6hTKA0fiDoFPorp0VdaWkPc1h6kKOu5BKPIysThoxe
9d2Ax0hi0AXR3i1b8YvQSwl8UkUyQPQWZUBEvE4q3Pi6D2Bavq1maLsXYbSg8DH0tM1tphCl4rVQ
74IFDJIxqAX0jk7LUXoocOsv35P/4q0I2x9iRXM02UdeRfiytvb/3XNmoDJseiTQurL8xThSsfk9
a0aFKC76itZy4iLj99Uzc5sNJJy1l2KmrcORrH8Iw/fN0qCd9sY3b3eMTclnNhe3RSYx1FBOpk0M
AbCXgX6EAaoPg428c6dYbJhIQTR3/VygIKmwJILEMkyjn6wR8eSwkbiCu5FIbtuLzmFISkcMF5zk
cjBrk9O+s9VIrlNt81IQ/ptG6kfEiN28xbMEoUizIZihudS+6TVEHUlADXzUxaDmP470/N2RDUzx
jsgmSVemUllIQneZxPN6r2yFDqAUO41oGkZntNONXg8nMMh5zMQpbik2dylu6R81/yP70K+TFXkf
NWMHP+zVttY3mba88nYbg8fTsINnhuAeiI195J8puaCPoiGbcmSk//Hr7/NeXyQgxgtCX1sTcphY
TJYzO4lOnJCfDLXWYZndPeFsF21A1eRvnApuLaF/FZywfR6Qek8JwFNIHQ==
`protect end_protected
