`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Wgy4Eb7y2sykqXgoGWHZutIX05T9vNdA/Dh1ekvDxJE8I9er6gvq+rnOEP1FQW2Ypec1SpEARHCv
1ORPhcWSbQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GGdAgKmhnR88hhmj/n/L95BaIrcFnpwSmJwHJ5EffhXpbgPKtXzep9n8tSny3fESxX6SCfNKgWqJ
KAVY3kJiHmjEwhrMidXeaadEe/ixovAITufbHnqAKy9pXQazkqAOGG3qQ8XWkI8FbdvM9MCbZcVK
JKCrHiPJKJVn1GF/2ns=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hthVdWNpx2AjyHLBKVPIQ9kMoQ8NMhskzHu8ZUY35Sq4t7+QlJsI9sV84jIVW8+6I767OLeBRVh5
VqufQvVy+iyA6uRqPODJok+OtPK/mmUY3yVYSGN6hiPljmRarYa3D1uN3THwi2N+VlDRR5Bcpwgm
4wK4sHvvL+X220ptpy/ZHsaaUPmSGuUNBGZJPvAQIzkmtzbVGcbbYFTRNZdvJNV3fJ2eXxl4QaDe
AGDEfq4vCNoEToYQCkezKpYmaKt+fh2PFAJM45w5EFBb6NddueyslDNseUhLfaREZbTrMCqtnELk
4yMz/uSU4rE8d43FwaQAAr4CPxNObhnEDDcknA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DJSc/fao6FDsBtUPDXiaQuyb1sw6O5ZCmlKfPzZUjK2Y647UoJQATV71FKC21STqAjIjXHeUU78q
lF3MIOtuA9CPoFTThNClRBR1a0nh/5DTcWnDYoxMU4+EFbGz4n3OvwJmsdsbb/F0CpOOT+ZcoeMw
I5zVGEHeaaMNu+77s14=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dVE2kzZ6gZQfQqlL00C4jjVWEjQEjXpHZaTPg6CZ2BKNSQW3todvojvfMQCWFv/mKdIH9j7gbGVz
BzRU2o1F3tkJImf68C9oy27qopg2sUTsot4T3sIhNn0oXRxPLMtt0C/q1Dz4TJjVQefGmODjIJ1g
v0f49RLcXq/d4OjSrYQn9y1UDIPnhy08Msw9XNqrt0xLF4d2C00mH/F3q6oo2ufdwMVuNp1W4vMK
HcpaXbQK8cPnkqjmCwkECVMGmQZVcECos4cZRTmmE34y6dKclBdMFj7/aU2Y/WJes0mvUSksUkLb
0PbkM88Y/IqG3+0XHLZ0cQ2IxY0bX0ppYag8Zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16592)
`protect data_block
UqSOjNseaHoXTt+Aktx8BcWVj1Hh+2xMMu1ydASnFk1PFtso+L+czefWICunV+WJYqQQQlHettcB
HFV4zIt05HezaWEWnJ1FmYQKSw0GqBonc5E2SjqiyJ5pPBKYJegM42xTjEa6GeQM2W3R8zJjdOlm
xMvq5zGq+fOeZvbvjnc7t1YH/VLvw52t+WsxXf0PvzfGe0CDBYbtadFL0i/dZnBmSC4G+21jQaFE
ndJTqSVoGODkh6vUDuTf0k4zksbz3G2uVTGqHWkt8C4CFMK4UW9kU0y5dVE/InA/hheswqquBUiy
QBdVl2UUk7ZI1qHvpXyptle7lOxKx+LkX0gV1/PzY2LI7bzceueIjiFbNexq/KcPi/FxVXmBa6r7
JcLO1XBS+0ZpW6RV481zGFqhDkO8FVZlGCeGdUgzyBDVvrN00wX8qwbS9UT9dS7Rh4Lm+SktI47f
yCLx9f6KTqzC+4hGyJWrr4v7opPG2GMgGahzU8ynefidaGJDEqxNYHXUfbpGO/CoHd8uFfVR375u
ljB+fWeY3eINh36O0QR8UqhLb0//zXjXB4bJYsaXzvoAuGjeYoX6x71FfLeaZmCQVbUnWV5qcdoZ
8VMmaoZ7bc1sgDaoJFmkUjKew+vqsg97l8JjRGA4c4rwXqOjQnsiHrHiBIdNi3u6NSYbLfebrD4s
46bbuHprtqYZuAY/ZXnVO/anZEAUhSfX049EU3KP5IO0nE0p3O41M1ho53oYidtHsQjQY3Mrh0q8
z4mP7pHOyTLXYrxAPtBcPVP2EMngFVylB8dyJG+JBv4hGmKFupRG+exwsekjThMEHoICRvQ11y5M
4UJLOM1rmcxFL4Xoi78iRlS0uvIuGnD7gpYuhF/IBYmuUWE6PAEweg4RmbKRiWeBnTjhdzCc3nGE
zdiPQ5QCNOgjx59klaDd9Shpw/ExlCs9t2Z8gEnw8xpSC/PXwfO7ySCXOD9pAQt64jQR5jXbAIu6
rOXAIFDfIboT48Z9qye/MpjDZkOyz2jNn2U3c7I5e55k6jh+9AUPooDY24kBe0/9eZcEIXzDATxh
MTikAWohHDq6BwMLr2TlAV7Uf2AvIDx+i3l6uWBFWmEb8SK9/WwP8T+NzHUs1Y9FlRLif2+T1Dog
MTnwYFJEQ9Ai5mb/ZwWgroR2uOawQmZT47Xxc6n0PBi6RExCcxjKNTYQZmkYeHmss54LGAjqVbFg
eIlwa/DZ5yA1H2T4imlvYjVKUVb/t8Ph3P72+igN/bXIzQAFWu90IBjKXBMrqGQG2QVIKJnNC+r7
frMU5OtyQxw6A+Ib+N/Uqn64gkI5uF5MDF8Nl1bO6g5O4URA6loLkK1YPMpbXwe3gpEZpi/zQgg0
6D27BCEggfAbcN4iSYyeunAluHp02Qnyjt2HaRgfCzcZ2g8uQVHyfcBv4o2z+TBulL8w7294jdna
trsgpkROmmY1d4Kb2toy4h3urfxtW8gU+HPr44L4x50h7eb26l/Tqo0SnkbLtELy7yXwpUvgd+A2
6kxteQfofhUjR429DdBmgNk8/E6EwRdBVY3aJ7ZsDRmU5PTuuqsUYHs6n1DP5gcUtxAKuSCGfsdT
SwMt6soX5QSYK0oBxoMADsKYis2PYKBoTU2mxmKr931jShps1XgeEi0BLToVhJ1+wJ1IIRYg9YQI
WSX+OZxAFoSAiioKdr/LbV7hTnnvtL/EXtlvZpuwDSLc2a50kV/EvPOkDwqfRVihm9McwZ1Uz06K
JdixWeASOuYTO8ZBgorGAR32uSPV4LTkO+ngRL4Yfnm9BScNglf/P7hSmR3qdSZL2+3V81oU1Q3n
4mP8gktgzFxQVVPyuyt5jxxyK9mXWNByUugYYuq2XoSJdX3D17YEpPZweXrwyK1ChvJfBzzzrG3K
68XCIX5eTQSGmFBNY2VCBbJCOTwK6yzSSbkTGIWRbe6/oHfuQsQKL9Hh7ir9KYSJcRGGeeDe7cco
wam988qrxg1mGvTcv8MK9dZPa4K4rjeEUMabBsA7MQ19QXHZdDopKoZQFsmDF9HVxfr5U425DDkp
RN8A837sqmPJdLz+QaK9W0hkNY3nto4lRhwhw9gk0jDiFsKTFC3AEkBkynLaH++gFGeAVOR4j7lS
MiV7ouRiPgOLci11bSoQxAR2PRprMKdKD/hQQ/HjLOIlO0Hn2+SEP5dswhc1FdF12BWbX3rzzrVV
L8/bzYxFYjth+uVRkJlWFecSz4oMgdlp5POum71uZCS3JWNl5SX2Jfee3xpBJUtEkQKWG1LQ8z6R
H8Q94dQ+4slyJd+IZdx5aTzyjiJxn+Ec7F8+UeevKeoApC04bJNv1hpOO/LDWS/PQ2PvenNabJ0M
Usn+5IC0NdgdR1M35LS+2GA0VVuQskxCMoKUkW+3r/pbXtM/bP3gXyIHE+9TBm9MXRbFGsY7Q4pY
rNME9AAMP/7fr8K8s5ALdjDHREH/e68I4MqVRB+lJoJ4ymPpc48oDpfG/HnL9OyjMsqZIRMRAcYW
Ebp+JJgC/6zeVq5bYDCaRk9DBhRx84SUzxygNZA1GMJcsIF3EWK2C8Mi/6DJOF/oFt94N3ZTWEba
elqSObVxFc5UU7KeswqLias2RsP0+wegOdSdrb+1brMrDeuwSIpciXt5hsRQhe/8+rRS6Wf8ADBw
AJCc3oGZxs2xVCkA7Z0aw/bZiJC/xVzwI8gHWIlnwScVbSRM6SAwADNk3eAeLKLCR2R7+dNOSiyo
G1/P4AeYDd+LWsaXubNWl5erLGF9wL7ex916NY9U/zO9QhqRuVmx36KiDllg0HistI2fQPvT3xMv
C8ttgYuq2EtNPv5JQps7vT19pTg1pcWtn8tgH1+WppIgEeFWgPjqSIR/7nRttMlM1F07VPKGW1HA
ZLQj6VFmtMegJb2jkxqsHEoG2INtEgrpu4TU6uuwO88fP6ssQiepAyyYy3H8v86Ggbx7i8PbjnCr
HJltqq/TkNp9fY6zN9Sq6oeVoJmjsRNxH4ltRsQ0/6YBiiEaEmQ4qUNaQlgXFXea15//LQQemsFh
uAb50281mOGMsHeWO5bmV4CRIjOLMNJZ4KMOepzrfz1U1G4LGir7SHAIgU9BsdVczbmrOc4A24z4
z14O89G6UfUvJbBLTd1HDxXY94xaL06DwuTfMZwSCFZyTZAJQOOR9GP1C6diSYTzK7fxVTQrZYsC
MXhWJyLjDjrqX7DB0wd06EdtNBGnf1KdSshS4Tb/FBxbqFF3kvKX4zYLo0rbX25as4MbXK5jRKYh
c2sNivHuiaBkNQKzFvCl7Dh1qy87tMQVt4FnWqt84uwysTNbdBBOdvShhc1cq3Ir0XJb8HCzK5OC
6UokLwuSfSt67/XHH3CSaVCltfrdP6STZSLG8cNw/g9oyvVkBiwvaxVGhxJINrSwF50fUOpsBNgb
c3As09inPQSQaDqMvXykmxlrCO1KHwLWA9fwfrexXGdkrc+IhIysSc+vRqTNc8soEKRX7OIIpMvc
EGcZ4AiETP2L9Z3ituTRZiUj/gggwEfiYwP8BOA0jkJElDEJaL2Nfa8TPsXR79uJq3prDVxMkeDH
XX2l+JTdTFVE/YjrbvAXF8ZgeyH4EMhYxGNXj1o2Ht1aZ828E6soP2kLd2iK/d9hFsdaFr2Xmh4h
zEGof5aEOxxXsNVJdYKSpALEy69kgtK+Pm5yeguKmLA1TpaRUZ+r7YCxHI7NbaV/trDRgz6UTyMp
WyKoo+Nv11rKgpgP7XeEjG1N3W7ybIxBNFiDKPgtlfQG4nnbFdcPb0vOv5vTyadnpIJbD7klVyAY
udinhBY205dtuMXqFvDmYCLfGXKGYIhDZhaDY/DuCuq8Zh06wmkQqcR3luhWtb9vKYFV5nXTJeX6
HwVH8ff0ncyTKmS58l5/SPqZwgnqsbEGS1Yfu3H1ahNB8WlGELxDe4dn7TzUQADbF9kfEd+MuDn2
18QSd+8vNpZ35dEEFuCaVDzJFB/GfC11wjybu66oAzCg1tRqgi+Ta0FTbkluG5ZVsDJQqodUzfWS
/hTKQdIDyDYPgjm40Kt9TThiu/IDyK3obTJfnVsg+zlsUjGygAYbJavKQJ3qwJ0xy7wNPMHr+8rO
3AnWxPRBHuQOjD3W6cuE/7NQaykD1Yc+df5TJ3KqhioOrO+eRj0J52vZDk4AyjpR8SmnCLUpu2iq
GXxcsf38oN1oapex26QKCVsQ+dZvtpQivbWN3EQ+sutZsojkdfii3vQZ4BPEL42gimf61JjJzyaO
cjPkd4Vv/2ILR78/jeiPKruMZpSbesfZ0E3hbxsu29FpmvHJwZJhYAZcds9VdadnxoAx4vs6Ynug
olZe5ZFx9TgmjPZ7HK5Idl0ZYw7DGYABEygVbo2ZW4f4rp0diod9h/GBqfjU6qwrNYlGr+BaKYLu
8leedtdQkXqD8FSUM+FXE21eXv3YKQ5Zg1T6JWbbVsnixq/3JIA9IYjzgQ3srwqUhuYEmxHt+7ck
CABIg/o5WliFRThzdf8zdVYdg6nf7bMEKp1VSuJC69iESQjPobVQI01RCP1JkC//6Pq1J/Dwv7/6
vCid/mV7MN8/t4uBFUrZ6JjvBRTAlPm0Om2BaHWI00XohPR34WF3r1TWEPRMm1Dv+gsbqqon5IrU
FKTqns63NzRKvrWO2xEP47kJi4/eZgKDKaXbKeIkpjzkpALf/d3cKZL4sdietJKYv5xvnOwmAvXo
HDgDoo+RVuMFNVd9nCkpA+x4me7cnENiL1v74joAGSybuNR/lWINTBfRa4H5ZFDQoKT4lRdvLVrL
1ZAQCNK76mQR3gM3Q7TUuSwYhkcp9y1mDKC40rkF79NOo3hPo/9ay+BNKaWKAKwskJLDJKy8WOsq
tn5VpsCDmTB3yTH4N9/Jm5+FAPPI27sSyj99zsx6f/4XR9k6Gk8quFQhFaDF3pZ+NnNF/UHUz7rA
qzBv105VWMWDvok+PaJHx/QYhCFDC9Gmv8PFiUJtMTIfJtcmuaQnPOE/gVDNO+iOSLpN7pZlGnBk
l2k1tJ2XGdxc14nMJJhbs64zQMg3b+06bQgw4WlWlfoDwuTY8insI0PLX8fMyTLAU8Fnq+lA7Pu7
8pdhwRYiXa5QvK9RWyXoWEPF/oi1TZYnCC6MgoA1cfnOBoxPua8J0uGtc3isIMO2Ah3VpV5XkwlF
+KWGX3oFdSP67xzGtEzoOr2sMqilfOOB6YvzAsI1i7MrjuOhUc7U8B+RAWXALoWGiBm1Hh/H9h2j
Znl+wt9AF5GtpPlP7FKcIou9rrVGIWjqe28aapfQoEM5qxfqi4LUly+xUBnBiiifCI95ey6nbF7z
rTMZJU+/yn8EChBOK1CaF/ntWXCUEKdmTfxHwp2VfuD2yqLmQ3ouTXwSX4M+U5p9OO486grRPdDp
3NRskG5RNUD0LtjEXDeibpjsL2DKVVo7k9xkgozCQM+39aNtWBK0zoBdSmqjvefmfVF6so2o32A3
HW+nkVlmPglZcroLzxaf/MjVIf2aRKsi2TU1I1AGnKm/cAmyXjiPR9VCBUqW26fG63Mo0728wr42
ebybQ2YYXmislwPklsoLoCVXU0XME2Dj3U9FlAlxQOT8M67VAGSD469tnKDFYSMehAgpC6bZhaGQ
YZIH5l/9dniO1wyjit/mmNj7JhHGBF39c239H1cDQ622mhgeB5bHEuDCC+6KRQCFhhQsWB+tqHfH
7d81Vsqoy/dUhxa/Wm7wIRBd+Z2agloAeXV45EPf8aJJTtw61zUTf2u2+q9uVVztdFh+NQgKbq/z
03XVbSw5QbpsLuOF/pRycmAUIqOmGnypYhEE2jch2L6XHbVZMRwXt5WvHbm1ydLOTLWmAnu4X7S1
uRoYsxjTo3r6p4kQo7Stg5mfc6pNYcyfU2d7D27oGa2qRJaFFGEm/wGJCvR55p8eO1DGgvin9KO2
4TifYnn0SVl+y4Fx88gS+pfELGGwHaa15Tb3Crq7hW6kv7Hq3ChsIzEc7rrWjy21bBKnXNrKv9yk
pggj3WTBSBvK0j4o2RXnPwcyjfUjjFT/1tyE/Ua39pOgMedaMja1frefud4OZwGc8Rnnw89NO5kP
OzzXVZilrAb3Ruq9uOBmXUwLX/cvmBGELmxcL4FdgVh4FFXsqzPoJ//zAt6UCBE++mDO0zg1oUag
DnA+baCecfKST6ZcEV1voaeqB3UNhPfcr/Jc/V+PvcpcqKAY/yYZRHNCttMAWSsfKu+zKBdpBa4/
dXPfJ1j6e7p20qillrQAjx8RocPQS4XgcXgKlU6lW1pTU6r/cqDIbDxIir0gixH1RYt6RPYj9Fjq
eRWrqkbqw+QNZIBQ6VLrSIecZfFpFVX1FLBiLfTVrq6xqHiki/lp6QhrvAQaFu8vuIdbPZx+SnvF
QeaL/L7L/gAnzD75nySAjwUF6Fvg/EhBRxSxvYectdjaKvFZpzPeWOvmZSfivlTMt+lTBu7JpzJ5
c5xBRU1J5DFlRqAIFLqK+NHgGAwUNQ2ffJeU4Enox3T8nhUYFjZxeaDP5g+ezEYU86AEC1HbMBta
bNJStg57fdA17f9HL+aW0jOI4VU1icoTlI8ELvnyjR0f2Gt/3QcYhB1XU7zIC2+TSqKUqhI/7TzF
OLtSKE8cpp5np2yLY7tp97X0CBROekt89OXGo8HQ4T5Z5xJVYO5jX9BvPBgGLxT3VLcGe6YaNNIe
Sufg/oawwvGv37qZgYRYD3Up4g30XCrz6wlDi9rstC9m4lIPSWfQaFSlbsqSXcRXPaJ+KIy5mMh0
CDSdgCIJ7BJCpbXZe2JzwpBZR8Zt5ZO4na9V2EMWrDP27aBqDldnNYhIWHeN4nygCMBQQTcUhnL8
s67aGd0E77GWN6TJCuc5NnQX15VwkoHfhrwZSCgm/0s1LmNiWi+95FTUzjLv6X6tD42Wgufhreaq
7Pan/FPbMaPRMS155qsOdmlDlgKDQKef/vz4lr/efEsI7vEvRH9gmQY3xUPJbSYjVK18kTP5+Sw8
29i1XOgLd9ESWxO+9AiFnSHwlbiJm9aT6WDtVi3w6EfFYc+i2SffQlG5y6A50y1LiwT3prDrK7CS
wDKR5zctPIGMzV7U/7jV6LJ/gGw7bVebSMRq8XClKutAfrdgGxKe2a/cUp6mDV2pRFCMXa+Lqb7/
KT3ouwMgMyBmAYxHJNONbQIw6945729iu9LtoHLvRnAGXVPIZyDGvG4q1/XpbmlcENKd6WaUPafA
zfrIygX0Wq6AcFAK48TUxdTubshb2jM/cP7WpLS/kxijL04yi95tP6bq2Dl7It8VQn/NUZiv1Sak
+LCX84JfrhTHCujzZxQ3IXoq7w1oV0HuIMQDlLlr3CzcZW000iNb+FYwNfx6NeNxe9M6WXSWorPy
5//bpX3tB7jh0HW9FHWvJAsRVEFEkhJl59WxxpzNPjxec4fFw7RjKMROxW0fSWt/OOWYfkrEhIzP
mRq5sYxkBqCYse0Z4AnUlwvlbLpB74t21BkS2XQwQM+cFsWGl0g89BlM8QOSfienEtZ/txScotHL
Vnxo0JPdtnKlQqbPrCqP3YA35zDJH371PQZjLBrTo7vWuK4TsViHt/XxZQCU97aE0KOBd9uliO4d
ZZO7jsmqVxn6m00bSKcg7WDzUuJsy5KSFnyb7ZsYuXGB7jTegat8pzvzaXfHLFvKn5/MMRf1DSZ9
JMeR+T0St2X5GkQAs3XFumg7TIo0kSbw41Cj1jRkY41R9p+bx//Qv542ncvkzrKkgdrIdaPCo9aR
SA0KBUHxF2MdDkE5X4P/51qVgzLpk9k6+tWGDeIPNhDdipzd1HQAYreFWTadg/bj2Nu5qRv6s8hT
Q/FEnL1wUNrdffzqgSv5Q9zZuZxsydEK91ZR8F25xNxOgDrzscx0nyalpvWgnv9CNLn+UX9R3Rkg
lvl2VVitTbGlhJpJD7rhnqM3Cc2/KP3hJIqcz652qyECw+HwkkUPbdsKE4gi6P53wpnBKhvoqdM/
X+CPAuW6x67eBaqV2Fhi6GRRKHEjNtqB2dFeOgtbVeLBn6ne/9ns90emBaabxyfXq1WnD85hy7Dd
bAtZkAiKzUKBvrU3TM9lRVmMH1bjBvEnTiW2I6OWH8a9SwdsXa5Nds2cozZCsRDqiGXJo7PR2AU0
sGhvWENGW0QPXE76IHdkjK7uMy9Zk8n5a3SvLSUIKqGLULWQYadx/vcQvAhYxbNxQcdOWSGSA6wT
XR6tUKtjhWU0pYdQoEkxaS0vdBzwi5r72qQJAksygLIu7IxSgQvmsL1T19LT9jMfyaI8dZU5mgX/
NQTV8J3YoXvZYdZ8GUyBTVmyYJFBi3EIjqqt3pII954rVeCWI16G/Q3LuSN7F3xFVfsG0lNiWD4A
Kusf9LPMJ4gSr/eYbg812LMDEhdTYtRmbpiZkxPY05kw6XJdoJ94vOjXvdlOt7HCr1105CM6YlBU
6UavV69HczlGjOQsnvzkQzctvUQNCMDKuKmn4oRCYgkg4iarVwzuCw52bpvIRtg/FMMinXPyZ+a9
Gu+KhrmkpS9HtPPY4T22NDMLkO77bIDr+6yge0/GCHZcjnXcgXQ5MdGBpM1hES2seidFqJeswGoS
Fn6RLmL1oPT5Doq5mVn25pEUPevzlAK/ss02yPYD9X48rGJW8qkoOH+pqd7+DO1mseg0mQWAm85P
zxWm9LN0LNGFtAOO1Y6DkVrT7aPIeDpcRBzZNlu8Ie0c83ybSgWVo2bXt+/sP0UKAnstN9sv1Kip
YWdLyTRfDSc2dXcbtT6AZ5fI1B5QlHxmWJyzwC0lN6gBSPOGn0vf5cQuEP/UIE6k6Cdg9h+ugD0l
qZHbebbTI/B20NTsTqIZ91ELOU7mScNB8k+xxtCMpFdc42K2ZdJpewo1V2EAIDNXam0EOqRD9AA0
Pw+ZuG8jiCPFAoJld1gSBbqvOGDjbyqPiP85dgCHJf38FiweuOr6xlNpfn0/10+2Sw9of3JosKum
ciEuhgQDyVGH7GjJOaoW8j34FF/r62u64B/ykPvc9NGJME4/7+0vlA0T6HWzhG7EBhtbABuBqjzi
gETCt0rP+YEemLyHX7EaP143qrng9DlQV0PwpMcKPxH/2qyxcC4v/cD5DGdKF2LrQdGwAzLFCIz4
n6b6E/N+WpplTZIatqvepGuvRPGbbIZuKRxOfMtvzjZfIwlTNgB8eftasIGxesPaBKyW8M3XsR/i
Af46V7yOKPl7uCuPAMdZ9pf3ZDECwnStoFC7kMFNnbZW5HC9SPsxWx0SaJfvMeCkdCib+aA6gfwv
CyZTnspNtOo7HPzSFcDo03ckTZwGpjW5GPYWiSMm2oVEHHixaPxZYITg24zrcOKgHGEjwfdexQVh
26cft49lk+GQk28rfDDaWsQpJwCZaKQdyGxBh75CCu1UdrCquk2oI5M/bglcPBedUDk4pk65/jho
eJclDr+o1NKcRhn+dfL23imxLUmzmT4IlYkvfJG8BiUYKTyZ6r6L/YCcBFZjy+Gs/ftFJXkaXijE
h+GmcMJLafP0D1XfpWyqVUrXnw3lSJF+oHLN5xkEJpj8EABkUaIttZTHzFOf/sFonU/dT9XFaKMz
ET9SvHoDW9d3deOwpK0I2yAkAmkkzkrvxDwYgq/rLzK9cknstgpuI8es9mSqNDqrIVM4tXQ0HYLQ
n3h6bzo3x40kmMVfTAA8snQUGR4vhzhdCbbOxhUdMJvmL0f4kM2ortXZsUL5HccFuGTZUP3V+i9w
/X1HnFIdsPBR/A73VJvy+v3HQcVcbHahWCUFp7vZSDxVIiPmNYMcvsntN02veGcFafvBpYZG4FBr
4Z8/Ks8V1lvxPrFxMUzM6eG/5w9CGabM600pJw2sjgXbIWd4FoKBV9dDP7+4ExuNhtN323i4TcYg
/cjCsMugWEZX6luZWOb0xI3QX0raUy7FcpfBrkjl2MfACeUSR+g6yQ0QgCLirX/43yTO0ZPVUSA2
+QXkyiKgBh54sp2zPjF6j5AnUa5tsNTqz4cCJyRZSWS3jB2KSiTpBXFrX0zdKOG0wNMhI+G4PMPm
59E8quCHR20iV6HZhBhfR8tnuRxHGeW0bBcrDnGCQMGKCBS1A0yef6hZfIgnomtTQrop5XK2GZbB
q/SRid3R1tPmRIPyfhqOOeEYwXqlj2tGrR2mX4fppC5NXSOJ20Q7JAUVyCfKV1FcRmxAFdYJ/nH9
MewtuVzhcBtrNfpfe06owd2Rynot+znL9xVkAV9eRy5sTvKcbLlRsQT5h/J/AZlXtUQi1YXcROJR
60xgcJ/Z4+gJWPyT9XP65ZQymloZDLAfqTpXIrnb43Z1gjPkg9Us3ihe0lu55ogM8B65vVIkS3cb
Zz++DNwf9S0PQ9wHMtEK3Kx4lE2dFKMaV4Mupuqvys/8Z8aRebd0WvAr4cJ2CQVkOsXfLYl9BMZ/
3OgCryts74NNWRdpgnsvE+xTiAXa7trjqg7elrI2jCdIqTMxtRnCfsatSlyPnuMCKsx4zxRDr/9h
w91d09WQYB04jqLTzeK+45cqUUO4aHYE7vC7jsmr6tD3eY3tcmAJUp8BzT4cOu1tcIli3pHreNOv
ZkKv9PkvX+3RxT4OAB8K2OczUHjal8oNux8N2dMtjZyQkhN1s+Lp4mA7CVdWbbMJzdV1gLNi/V57
XkmI9vFg106QXmpB5vEF0hQ0XDdm/uRvtBndZ8XLbGXIm/Q/Wz9niMI6uVAvnO4Z6vGJHWEZuVGd
2+31NR7zQJRsi5XPcIUqQjWRtQ19OGUcPAWf/nijBRNblMUvE+NSJ2GywmAW8ovpMRstjyW+Gowd
amxuv9BcFJRz/0QWDlFv6CGQknalzLKSayubekhJoJFWt2gMlzwqgeWC3mhmRGZjvJKGOwinvtgB
DpSPEU8Gzo48H9IcaYirj7JF+lN+G+LzHLLLZPCoOJA5+OeUM+QkaFuMwNXHfY1KWrj+Rbn+iDiT
yBhpWzvFIUIzk3RJlknA+Z0tAMjYybqFs8zwTQk4v6rcAuFy3m9ePYSYKbmfOqInaoDfJrV9aUrP
5w4rRbci71W3K5XCPSEz6aNMIwOCmA2ExAFfc1Q66Nvyp4CbwBWLDo2MDqr+cPu2AquANwQ5E+YG
1pK+2nCBEanr7JqmmN1vsHuLP7zboGYxg/Xg6uvUPvLJ1gRRxQxg7hHchaOpF1tWnWkZ41F/46zN
LHE52kaWNGZC/m9P/R06sM1jYPoYgUBQRbaDz0YUNlfNpKku02MUPS3+qhYcoUkhG3axieXNAVaD
NoiXCEmEjnAuAbcZeGOHJI3rDlAJlQRfyqYH1gfJvJz1nJZMgEuCbIRJ5QPCbdHUvTeZhZpaWig3
ivy4pIIG4W90snER1MSWtxV4U9Z0CdpEJRw33t+cU+7yd823poHzgM+L0/YIkqSQBwPjDtSskIEP
fkUFa+IvSspa+DM08cShPyzqkeJlLWBcGzxtnrAlG55bvKKt1C6M87/bkyySR6bSMdvbjUem0ins
bUn1nltIPwMnnMmvv7wGOi9CMafaTIwPzSOqlTznL/co2HzdR8wxsXtEQB+q01kizSJ/KmsdmE6B
5j1pQUko3b1Smvoj+jPA6veZD4KevTMF2S2mS2rf/YCiOYzxp3YnBkLC5KOb76CVzlFfv2M5oMX/
QQnkZdr6mmvE+V3Z9wzCMsMLo5c2m6uRWxo8atHAV4su/MAz4p3tJqeN60U6GzOvODMzIK717uCT
Yrq7AScZm2WSYxeIkRBuKkh85+szCvcLm9nZz2T3Dfm3AW4crlHw0e8aCXAfabdxz5NAZBICSd3A
85AX5Fx9QRmpybVkmZuufdjbaB2Ul25Xs6dyyJIdB5syXVdV1pLHyDfjPgOffzOo7q1U0PCC6K8+
OMJz0mFdOaOJHsHyj8u5xMMRDq+si2zkB6Z5hoS6wfY43SES83xJCCJSujOMER16PzG5z2IRFbTY
v7Tx/aAS7v2oh3awdkkef8HIQ/OrUdysZOmxJXjq5+YHd8qNS2hRiYrmHVzNrphgb7pfJXvaqFk4
gPr2Q0Goz7u44PZ/18zJG8DAcby881w3PB6pktTrjGyIoZgsHA1QaUpMhPBKzo52mRgeYmJlpmOn
2bAUuNiauzxSMfNzqJjqfMBKz+dQ5yrJNqKFgo2t/kphhEVADtFJwlx4IC4lMKjI/pAt0nuj+QZb
B5AlTfsWCNlalp78UTSpicJcmMxtWfFoK5l1DeZu3pOKkqTGuSHZJF9O59OZ3DJdRMpLQmg+zaPz
3czZPjTuvGLbxa5IfBT6LmFC9aox73YqmDVJhUHIsLy6TZlgpkRE83LpYPCkfhkUoep/L3u2eoGs
PXLiZF3Unf+nuwjj7NkSTQlJ/+grwqGkJ+GCEwJAokHqn7dNOfcSKWtTqdoRRg8UKlzw80HqVcFK
6H6cYTaxEEVoniE5nO+UThz+0Wku6WgVzJHy/2xqWJAsPqSSPhoytbwFCkaAMXKpRM8PQ0Od65kH
0+za4TPr6xL/yudGYczrwRCA4GWix3y50fdQZbCyuaIguIdewvMCmmzXc1sfIdB39cedoe4dkuos
u94Q6sntMh1P9HQmogwD/lm4wU4qv0+9BMnzbOK1UapoxE5KvViYmZhOjrci9+KqwBpiLJClQxFJ
gEeF2sn0LmhcKF0XDJmMKikf4NVuMfDhOYgkWrIQdSQG5JDyxODz2CQqq4+TGlJIvPQeeWNdRmFu
8RLfGcUFxYEfTMqNraDzEfZlPOFV8/XFtf+LNxg6UF9CxGUizixq22WTRAFp6QFiSVcfgrdr24yI
r2Q50+dx289VViR8mva5R4sUb3iq72tX1IzPO6ZqfIrng7cF1vCwbRvE4e6mYQkBemNLdEh7a007
Ii485HYcXDmQVkzDnl1C452qfvrll/9ViNNwa8n1i7Q9oQdl5C8kgcV3xlfUF+JFq1aqi+COUh2P
KL6IVtVl3zdEg1NXmb8EmU5/Jpa+aKxjk8xqS1oNNvM2vwhuTpNW5U6MamFshtHHqnx2LoxHTdFD
Yno2PiD0SGnT8vFscghh/gj8dZpqJxtO7nYSCK4uoeKQXYlYmcRLH581y/5BlVRZ84WpZmMAXKDW
cYPNpRDqytf31qT7H40HWBi0fOi7VgEFLqps7+9154HLTIb6KG837WE4HrLKuEpr89B++hw9djlC
yojMkoUgWaD0AHECOx6WkVFQpkTVbM9Cygt830DXsdc4xwEy5i22ST/ukfHWH0DOLHG1tA3GBlK/
UbmSRvVc9/aHyLKE6FzGHqtaFJr06/JF2yO3FOSedRzNGHx7XEetAQJFB28ayKUYBKfN2cgGU4NW
FReYFOjNGie7QJ79FUx0Ws9YZdKU4lW0Cr8NymQd6JDTYhDuQ0T5x178XInHgYQCMVX6TpAwib8f
dUtiqvwXKih1I1C9k8bGL528SqIxc6Y+xvVAA5m2Ja35ak53R8wePIiiuVgQm9MfiWK/bxHkj5zI
K+PkodwkQ5QTeWR56sZ8Re2rzTLFGP8zss6wpikhLffJ6WZ2HT1jhYp9eZPj/TLHQrBGvOChiFGd
Y7Ea/1UskX6jbOMFTkl+VA+lJXMmDQrMU/hyYrd/2AEBMxkq3gn9tVgeJxmEuv7RgBiF7XNazais
L7I7uNfq9guQqHkdCiUt4K2r+t3v01cYK63GqVj1LIs0kfFr6hF6XBcI/8qUMjUGsnZpsZ7ACsOQ
bPTzwIOxkkCe/TvX6Mu+5jdbGXNApDWxXCmA7cgiLv33NL3iSs/LLYg5XvxXwbpHFmyY5i2xFL8W
cm5k/+EejVW2/rLx2ON5PoQ+h8tokLJsjTKH3Px3kydWo6F1KhtTGDpHvkXEL5u4CDvzXv5RU3XE
scQ2UptPg/h2RxU5gocn7m6OZY1roqOIzLTPXT3nnuspKGOfwDDz+q7LaFcLZdbgEhtqZn1BuX2c
F9Q+7SGkVMhH28GEPofhp0Xq+c1Qjjn20XRAoeU772fY4pLpBgcGhmPuMCnHRCNV4a4V24J+AfdA
b/RXMobN+HOo3F79d6oQotOio4XVrDYDxJeKFU8xERC0ahbSLG4YlvffIbimHWhfpqIf0NT8vwKs
TbCa8F2QzAePLgZAKYHh6BFKQdOhePhWGWXzxMRSzIY2orsfSFNPtekq/qajx1qtMOY3L9P7VBPf
Jp6qZlnpH4KAW6TktFzMBoWdKKmHM5zQmu7EVWbwVHz/gUNMd7p6kzniyK7P019DaH2QmRm5N+CQ
DMkqBmsBP3U1nBrt7rhjlFLUlBJ0IK1gMrulSmYTXlTwpRH3noW5xMlF04A7ecdzX21jw3vohWoZ
ITtceSTxvz4gYbBTVu5nY7UwBEBdxYaFdrsFL71FIbQFOjb9Y5wgQXHsp8Q6JcuKCIaPDHfd9fWP
FfxT8RPSENbH8ubuzjl2kTTStkSMIXBg+cdPwu8K9TuOsSKvwKSdqY9qimF3DQ+ZLpgOdywaSnWz
OFRZWQ53AVf8xPDCuvaAAW2RNMJPDwEGcjU0Zc72WNYUuPFiUWGM/pRWRp+P47FLY3Fbr8CcyLa1
o//KJXuZiW1ZK5VVVve8EFbfg6u3VPbDoPGt6UUDz8Diok2qqHVsqvxuFXatcu7bLU0/BYpmFEOl
LNt1S24deF2pF3/eH2/Dmml9xJmzIV9kHwvJSqFb0Ta+DiD7iLgfoatGtzZ6ukGTRada0PlDz1Tt
y4srMLqqZm1KA5vHq4mW3JQezJ5LejnZenxLB0SaSZHBGPSG4KR9yHXTZ9SRo2wvnbcocpTc0KAt
rOK+4fiY353qLKUBvzsuiQ6KAhaX+X4ci4SyAjMyxps6x9M+bXDo4wXFLwnjsi7oaCe41CnDehii
W743UvrTgpoHUXlZY4nktMmrGUYROAxU9eaZ/d4/wyWtYo+BxdAogbK9vFNwjnvIay7MuW+ALO9d
DYUgFX++jm2xVsAR6PG5lAoqkIEwp1zgJXubXvvd3acpWbOyohTur0TYuu3/QSCUSiBGJt2kDTgs
pLFPUAvptc91RgM9Hth6cRCZ+WJ+3CUnoZxtGMXZ6PVYYpJYTpvH9yPdA/lMQuC+blmOJ7a3lIQd
9V3y7JVNroSokxD9MD1G/1CurTbTDTjAoaAhqgPn7chl38HNTExfPs8C6/JhEmzRNUxRePENZcCe
IV79CsuEf6LleuAgPav/vgOggeZpGgwsleuiu/Cca59uKMBCyiTk8wIUw54vqoO9o7aUq778DGMe
vfk8bMjWeNTMKOBfVm6cdHHsvhLVUPLkvCrqz+GRq9LdcTCHsngg9wVwOQHRNsv5dwpJnZblP/dP
w6TllR0pDEEI3563+Kuxe2hUeab+CFa3zX3QnAk74GegkzOmWbtT7gVICGblzokw+oZEOe9/6/G9
vkFWSCjmVsKWylkLl0RcNEVsSv853tB0u3nGKeSM2x8cXOcVMoZ0yqBvi8FvFEZDcksqqONXiv2Z
zN6X+wem/ECSZClyLCmm/KOOdPpjxzlhmAPNkMXdVJLOg18mBXOIKRkDFrDL5ciAuyoGAgkTWBbH
i8EZhlbmHIiEPuOAfRVR7MIOw01Bj5OgisHi7Xm39fEw1DZLfdSqzrtmIxnQX01gShRPReCMdrPb
lmEUM7gtw19Mvs/4yi2wgyifEISebJviRRmE08I1bwUGqUltCZoz3V29CTSsFD+gM/MXsKQwWhiK
cOiUrdozTAMQVWxmDji1DXG5b6TqTm0pxNymqzjZyqqxuppdkWH0SlDpmuT+CXEURMu47D4bVp93
YNdv4PxzHRl/NlxyEzub8s8B256RWsTeq1iO9zc9ayhkPXpc1hzTl6exzl/HOfQBtlyBKLH9NWJg
7sTYTGAI2t6Q303vbM+ZODH2scV7f9nMbh2W++NuSUCaMhG6mWzfvlf240C3M51G8GxG6QFIImOt
biGSwzDgXVhmd8byOW7Ctlz9aRq/FgMdNJIxfQiAhOL2rRawOdevfjuY20WDWReo7boRiAdJUCNG
zy4FSGZ5Gc/5PJ85WPtvY6HJGYxXOMh2D/F6F5h2d7gtg1VIeNV20jzhMZazXnZwEM0SYwzBSixH
jVUt6xq120xeunuHCPCDOuoZAmnPOLZ3FMXnMKdAxT0NZBiCmVFh9qb63qEzzThXd2i4Exe67gQ7
kVgodOF16mdwkzMJ/jbEXEN+WTnpSPuJE/+Jc32ZPJU008ASZ3kl41Vqy3BkTSz6RN+IwW7COpE2
6jcAHbsmb/dA2CGSxIr1511etao11m1KmU7KLegDCToEmxm8NtQ1tedcjBNibRUeRZvHRJT0KbRH
S83sgkC0wwojOwDMDHdUCddhUZchEwLqcD+KOTFddYgme4ClD85KzkjXTInNzqPNFPnjW6quqJbI
HxuBXOnRPsJ2HTUtPNheEomt3Hn0i81S8T/SP1qqFuh2x+ZG4d205HR3+fzEIpLmL2/DO4d+1xEh
y76lccBD2iXGSYJs40ULWWlDor2EOoRJZ8KaToKiIR3PQ1kY/oNxFeYIyVQ5kKrd99HhKT8j4aNq
FwTKeScZfS5knUrMp9JaKgboZZBkrWuqGbkWlxTG9sdxJG0YqCuY2cWQWr3cD8Dn2Rw83kA24S/n
Ex9ERuzNVGiNmSKR3OsIdXM88rP2yyyZIqjKntaD4Iom7ii1CTQAH/xoNvXV+Tt0aq+6xMRUQcDw
ajEeG5OeSfMiC7kmK+FCEHGtxdUodDNk4o41zeNG5i3vptClUDyvVzuH/aRFrNJpnz70207arD7n
igByJDIDGXG8VS3fwgCR9iRNeccpeUQwzO/U2JcY5x7eo5ATg01XoiHnYMjlHZW5nBxfVYKJmxRX
7WLyhrGBFr7bTbJfkKorLFix554e+ONXUJaw5dxXklGe9lH4s7ylqg73ClS8fd/SYsC5T0qJw24X
ndadxPUPihXCuMpWzwhh2MsTSzywqIDu6KrNJxra7iwbHrN/aMe2SPw7wNQ4AspvZ1UjlSP/6F/c
aaUTxcWZQi8kmszid6TYAU5OZd5qa2Swav4KkITuUVTnYxhYxpZGJWCSLUsX0NAK/Cq0hkKMIURJ
mm+nEfAVnHnSgl+e7SzqqnO4HaSuV9LmIY6YaPPwSmQApIlJT0TG7BNqmnbT3OGDGx4eU2/lFxng
TZiXo+e/Q6EzsFN4FT791qiQKZXDkQl+Ti8borptdjX6eo/2QnRK63EilQYa4aVQzOueasrXMLaP
1Dte4c3RTHIOqjLdVajlFtFJPUbKZIRxGVQrPl8aGEhXMq2DaRoOIw06yETpWiQrD62fhlhwCTr9
nLqL9WZDRcnkAZQJ0etwOWfMwb5itw5UDm2cYHobdRfvuEPpHa7kKEpapno8Y1EaXSusBw95SkAi
hCyv6QD3mUQSbduIU0bRxQf8OiVY1X8Ovgj8cjYXIzoICauxbPksIovaNjcpfgsDcSFs9qgXLHpz
aqNa3S7vuLoN0Oh1gFg+6JFEsk88NMts+uLaiR6w1xLLOHUMxr9E5zuAb4b9N0rI8gL0qKlfG4Mt
8qsiRmirXy9siEz7EGWroC4Ur45M/0Otg+uIJDYHwLWjbeFQ09nrLbWUeWondKiwlSlSfaXg4Bb3
D8ygZs07vcL8Iw8f9oM3r+0kU4QOf4WP3LD+idZB7El5kuHNnw3LF6elZcWOa2OUl/ZP0HD/DoLW
tIUjGFcuU3bI3mtUk2/d/XMOTJrO6Wv0qZhOaHdALuvefyxY4JuRBKp450DFCuh5VZWjwNUe0zPn
fIA5havqy9uUk5qtF1UC8dAoKjklOAogSXfta1voOz8uwgjpFsbe0ZAK7V+k+H/r/IargYnDtyOq
XG5d4EuPiuJHxdzgoWe/zrumhH9R3IgJN1Wpjnr7SACWPGoe03JgOPJGECWdhj1Uvnhnj4iJdPmc
TI0p/tB0Iy+Y9B6Ma/xIqNwCxFJpjfMyL1tBMMTRyep2CAoL+DdKzky1kvQBEo2hXRFYoxsN2SV0
/dSP4XV9wTnTyc7ebXXKUfb72iWKmF+r2TOj4Y/5y9sEVwQpynzENugCqDNM3wBKMv0+XvMuEIJ5
NcKBVUlK3pME259LFkskxVLjTQrlnlxd41yNN2Rg2JFGSHZCN3mq8ocphtT0vcnehqASKjR7B7Gv
Re/5/QRHZhpyF+k+PGORiUfnWF4YfdJ+DyBEHIl2YBaUQc6jVRo0HkQ450iV5Jy4lvJyxIYl5Mwm
n9ZaqjG5oHZIOOhNYfjLI89J5iLEb3EFtsAkDVnYRCdMivwlrUHQHRnQ3oDAN/W0o1+m65ohQ69u
ytQbsPyLLATbb9RdCvTljy0Np2NaME5T3z1x7Xq5ZV5gQM2UYRo9muSMxYq83mmIX1d3myfBnp+X
3pLknykv3YkQ6+YWMY10gC6Ls4BNu/2TvKfhHnQlMcpyhU3cDzWDwib+u34OzE5JSzzYVrALT3vL
qjtqYg9bYmuiozIjcPtSjqom5rq640Ju+TZa9Yzx7/y5cMlMqcz9xxw8BibE1AozakrVI0UHFn/j
ge8SBIWj1hYNlJsVDFBjdVL1Ah6mMRapQfbDJN7Ruo+fS0SbfjNrvVYbhGkKGWRh2hWwOQ6UQBsg
lP561UTwtpzDh0DVLgr8ypOkMOX/C46J+ZK2GCff7PYmJJHJPgL0A5OpbjkXKX1byqIKCUcPI8l/
MlY0cM65KwBDniixle7LbcHRDuedz9PLB6lqV8Spz7TIXp5JjLOF5mhnNnZqQ9evlIur4vzRRzbR
9ToX0BxyNDJuVMmEi2rK0D+LVAkwrhRJfX2Gksbiwv8XsAAQykqWXU0M0iZI6zwbQ2byac+4w6in
NE7BD7hgSY6Io4dy9prOCjXV0LKIXyRHhX2CAzvHKU2OcUMs0RRz32NN3f4as7nAoV4+7DLyJH0s
JU/9VGBzMpAJLSrneHe4qdFbylogCtKDmvjXyGoiqxBLROgmTvwwO1M2cUJmBMQVwvgFDKlylqUL
iXRgxfhpFGZn9VTIwUlBRVkrY3HGUrJ0yGbvchJzD5AEYlF3jB/42TzEVEv2kAJnXJhXCqDSsny+
P0FyyElg31/zfLjD/Ezog5X1ypelo9+Jtvc6DOJ2WiUWvFoCQYYyXy47jTYfTRf9M3rZCe2oy2bP
T0OLZ2EwJTxA4g9lQcVPZ9qG6ZHEowAKzmdIXeojIfz3caA2NgHaQcjnq6By+D0QlMOJxQY9CLGp
WSFyrS4jjhlb5meQ7VbT5YJQ65BeRvvCtpPJ3F1BN3JSXdA+Pi7RFIc1heo9Y8VGyCxUJKbeKZuj
q5zwz8p1ojz7bUOEDWZPzam7mt/i1TY1u7+HiKpQr8dCfJbA2QQe6X9JC6R4+Lwm10ZLLyhzP/dq
Rm1dmy3KbQZoNLj2qrNRx/ZNjw+1iGc1tbBP9U7ocPE6jyBc3q+qbEMq/g/iGkK4nm7Ys39Os66K
DOjz7wN1gCotyEnzLjc54ZBxRNJg5282iAeYOHNZUsIiH7guBBj/3LHVmUrAO0jQqpVfyaFuR3AJ
BVFwrZkUaTnQamZoWZqICjoPMuPOsWymWOHZCrnbuzCEpqXx2xaWpvvS7BP34fIEbPAkwu21Xc2F
9iRvBV/5KsOFjwtt3auNxPGUp+DHXnvRkd3sopnIfsPXCoKH9HsQYzgiugwWugdKiCzw5oaZBEDa
YYd10qMZ5unl8lMdZNPHA0hmmSMDPsjTrPAybMMRP6KgXRUNkt8N2UXezLZ5JK+D/3Wk74bs6L5s
4cuin316wqXUktO4sZObjiyuCCQGnHjmZ0lbvj7XcoZIVgIOYxGxAaUhsS0TsX3O8yl8rbQqe+i7
R/V13BR5k0UNY80jnKDBoZcMK1SSxrnUz83rEGs9TBFNk9kcWamD4t/LsLwt1zowrCNs632bDhpe
iBKGmf09JoY1e2J+GqwjhtAaK5kO+CwwXoffXlLGCsRUby6jAn/Henhcpi0TW9vooIbdARuWrIM2
kg3bKEj5LOKfqspH3ntPfYNfYZ1RPpcgf6NmpKJrAEtpN/l87N4eIS3Dxnfc9t/LQqCgZ4Ahn9/S
MLYki2AkT45A5CntQ7R4Eq0o5MZ9L/cvMIXZRoRP7ZbW0CiEcWQIwk8VD+X9lpjYSmKVZDmGks0S
eNBiCj8PVIeUJM+yGQhwklunGPlqNnVAd1CIOBTSPzcaSZka1e5j+MQKANRSXfX4WZzVGkOwv4oc
TbnmUhIt2SHnXMi3rzNXxXgk4bHdUzlq/8JpCoejM2/AijBGdm7TVD7PUKTnJz/i2CE/P59gBmC4
1NvAGM7rXdjyGWQaVBzZHAkc57YcBNbhBx01NCfECP+Um72rY2+/BeZNIw0v0LMSPiapAdSEo+nP
iWF4ymXWL78s+50hjYy851z5Why2reMxmMMr2jwa0A9af5eSwPGPqL/bai8SJGtMIgGgY6YH8UAm
Okqkakw7Rm8KFxaB8NVzZtXp60/XZCm+uAKu5S+Vq2DVw1edWSE/ioE9CSzyWt/u1V7Q5DwyHCEu
xcFiR0wBmuJr47z+p8ohYxwEpuhiRutM6GBlk1v7d5XGAGfUr/t4f1+CGtCfjBPxQTDuI16WVC7D
MdVcucWhe7DplYLXkShM4QRNgJsIkCAMRcVWoXg2OG+U41NeLDMUxN7Ci9UtOpSoNldWF0evIriP
3mrgJQJhFX1UQLY/XaUrcNuvVAhpKkbUjY3xMMviDn/Wr9/8HU/DEaHzyPqkn6BQxZmT0m15Y+3I
jACzzPohdrd8cUed8bT0L99w7qK0Z08nxJbMd9URKrkNfg2rJcgq4r4fHHOT9OUe5MRmQJEaTh3t
X7/STA23QyeI1F4k8XDlHFZbuMwFJlLVKgmzz739uC7gxgTBV8rMMp5iZg7QnlFp6tyvqM57NK/9
rTzUVgrg38gA36+3A+7yg/JOOci20dIfrpDV0PIz1tnl6avmhPuseOMmSk9ndzPMMEfej5XgeRVe
zmvWcFIhO9AslBK5pytoIorJfhWucCmr4JCsLzzs6yTfteQBp+HqlMVblGLdBGjNfc16DFygsPOq
dmNHOuzz+FDZ1NCe9hgFyILbAkRKeiYxD9Ql+FQIxJMUZo6zpqBL2kGK+liyHAw1FLXI5CPuusvt
k/7D74FkFzL6jcFvneOehXELg2OKaWQtIvCh0UID2k00jAWiVSFkDxNleDH3mXEXLK7w/atu3SzA
mfAu98Xb53lk+w6BdlTnzeH6cr8eyzpsGOmPP6ZpldHVzqSsg5XZxNt3YK2PUkTURcvbW6+rK9Vj
P44UXsh1FB5pBeckdkxaqCMY+pZ76gHMXHWVHHqRI4+M5n49iVuNieY6JhHFDMNLr2u2pGplfw4+
RpnYA4cFmB9F68tazb+E5296DyTEE3ziVsHXbJNJsD2BtbvM/Gt8X8z/TRXJbB9kDsYdmSQkXa0K
JoE3dEjolkLalmagUXRtAT/KwAllq4WxUH87s3odZueKNTLKsx6oIy/mKxI5lZdXA5QjEo+iFq96
zBH/g8zEMPzJXuG/5yLirynmmC2GiAjr2iwmSlfvscvqb0aFyxx/Vw3TxXBnmaiuZeks4EXlzNkG
74dickZHFC4HBtRTVNfQA4eVZvJi55Vt72KHAfWqIW5fBOkLwSPuHew4sBcWDaQULVgYffe+VrKN
kceMt+waxbvBpdtrphdC6GemGEomEdVoj97NGtwPJ8IKTf27haI9B0/hi8hpwFGjiSg54SP5X9w2
UFDKQ3NTuUtNvloNwsehJ4p1pYhcXFYYLCh1Lh28a627LY3T6LMt5qtrng+Is7leOZ9rD0Ect+i2
xgk5fJJelCMPUwwQNvtna2DVYyG8Op74tmDzi7pT2GWxkwcssE+chcIB7zSq4GknyDsQY6EwBkB+
CyuuJiK63YdAdQg39s/s7NQfbwY1Tov3JD9P+nr5WTK0SqdxIc6VKCpAzhfFr0Tcz6vrP93f9HVV
SyVUaD0GOOFSSZYhgkvysyzZZyeKtS0tw1sJfymyClZvgXLSgugEMSGyesCnd58QyJhEHgkqQD9w
ZK7SNQEksIXf7UvkMkPgzx/MxTxuoPIKJmDcRTuItaG8AqhmqtWKoKeNhCdvdx4vdq3dg/Ua+fXb
xhuhhCvYShCEVGhs+C4cP8vr0jU9Ic7hQF6MYMhPBJ84hUoAFLeBjsFPQSy/lPYlfVNw5AuxCNXu
TXCOiAk=
`protect end_protected
